magic
tech sky130A
magscale 1 2
timestamp 1528465711
<< checkpaint >>
rect -1140 -7670 12104 20989
<< via1 >>
rect 3735 12237 3787 12289
rect 3799 12237 3851 12289
rect 3863 12237 3915 12289
rect 3927 12237 3979 12289
rect 4103 12237 4155 12289
rect 4167 12237 4219 12289
rect 4231 12237 4283 12289
rect 4409 12236 4461 12288
rect 6469 12237 6521 12289
rect 6533 12237 6585 12289
rect 6597 12237 6649 12289
rect 6661 12237 6713 12289
rect 6837 12237 6889 12289
rect 6901 12237 6953 12289
rect 6965 12237 7017 12289
rect 7143 12236 7195 12288
rect 3735 12147 3787 12199
rect 3799 12147 3851 12199
rect 3863 12147 3915 12199
rect 3927 12147 3979 12199
rect 4103 12147 4155 12199
rect 4167 12147 4219 12199
rect 4231 12147 4283 12199
rect 4409 12146 4461 12198
rect 6469 12147 6521 12199
rect 6533 12147 6585 12199
rect 6597 12147 6649 12199
rect 6661 12147 6713 12199
rect 6837 12147 6889 12199
rect 6901 12147 6953 12199
rect 6965 12147 7017 12199
rect 7143 12146 7195 12198
<< metal2 >>
rect 5289 12607 5401 13913
rect 5933 12713 6045 13913
rect 5147 12579 5401 12607
rect 3723 12289 4480 12296
rect 3723 12237 3735 12289
rect 3787 12287 3799 12289
rect 3851 12287 3863 12289
rect 3915 12287 3927 12289
rect 3979 12287 4103 12289
rect 4155 12287 4167 12289
rect 4219 12287 4231 12289
rect 4283 12288 4480 12289
rect 4283 12287 4409 12288
rect 3794 12237 3799 12287
rect 4034 12237 4103 12287
rect 4160 12237 4167 12287
rect 3723 12231 3738 12237
rect 3794 12231 3818 12237
rect 3874 12231 3898 12237
rect 3954 12231 3978 12237
rect 4034 12231 4104 12237
rect 4160 12231 4184 12237
rect 4240 12231 4264 12237
rect 4320 12231 4344 12287
rect 4400 12236 4409 12287
rect 4461 12236 4480 12288
rect 4400 12231 4480 12236
rect 3723 12199 4480 12231
rect 3723 12147 3735 12199
rect 3787 12168 3799 12199
rect 3851 12168 3863 12199
rect 3915 12168 3927 12199
rect 3979 12168 4103 12199
rect 4155 12168 4167 12199
rect 4219 12168 4231 12199
rect 4283 12198 4480 12199
rect 4283 12168 4409 12198
rect 3794 12147 3799 12168
rect 4034 12147 4103 12168
rect 4160 12147 4167 12168
rect 3723 12112 3738 12147
rect 3794 12112 3818 12147
rect 3874 12112 3898 12147
rect 3954 12112 3978 12147
rect 4034 12112 4104 12147
rect 4160 12112 4184 12147
rect 4240 12112 4264 12147
rect 4320 12112 4344 12168
rect 4400 12146 4409 12168
rect 4461 12146 4480 12198
rect 5147 12170 5175 12579
rect 5289 12473 5401 12579
rect 5924 12473 6045 12713
rect 5924 12471 5952 12473
rect 5883 12443 5952 12471
rect 5883 12170 5911 12443
rect 6453 12289 7210 12296
rect 6453 12287 6469 12289
rect 6521 12287 6533 12289
rect 6585 12287 6597 12289
rect 6649 12287 6661 12289
rect 6713 12287 6837 12289
rect 6889 12287 6901 12289
rect 6953 12287 6965 12289
rect 7017 12288 7210 12289
rect 7017 12287 7143 12288
rect 6453 12231 6468 12287
rect 6524 12237 6533 12287
rect 6524 12231 6548 12237
rect 6604 12231 6628 12237
rect 6684 12231 6708 12237
rect 6764 12231 6834 12287
rect 6890 12237 6901 12287
rect 6890 12231 6914 12237
rect 6970 12231 6994 12237
rect 7050 12231 7074 12287
rect 7130 12236 7143 12287
rect 7195 12236 7210 12288
rect 7130 12231 7210 12236
rect 6453 12199 7210 12231
rect 4400 12112 4480 12146
rect 3723 12096 4480 12112
rect 6453 12168 6469 12199
rect 6521 12168 6533 12199
rect 6585 12168 6597 12199
rect 6649 12168 6661 12199
rect 6713 12168 6837 12199
rect 6889 12168 6901 12199
rect 6953 12168 6965 12199
rect 7017 12198 7210 12199
rect 7017 12168 7143 12198
rect 6453 12112 6468 12168
rect 6524 12147 6533 12168
rect 6524 12112 6548 12147
rect 6604 12112 6628 12147
rect 6684 12112 6708 12147
rect 6764 12112 6834 12168
rect 6890 12147 6901 12168
rect 6890 12112 6914 12147
rect 6970 12112 6994 12147
rect 7050 12112 7074 12168
rect 7130 12146 7143 12168
rect 7195 12146 7210 12198
rect 7130 12112 7210 12146
rect 6453 12096 7210 12112
<< via2 >>
rect 3738 12237 3787 12287
rect 3787 12237 3794 12287
rect 3818 12237 3851 12287
rect 3851 12237 3863 12287
rect 3863 12237 3874 12287
rect 3898 12237 3915 12287
rect 3915 12237 3927 12287
rect 3927 12237 3954 12287
rect 3978 12237 3979 12287
rect 3979 12237 4034 12287
rect 4104 12237 4155 12287
rect 4155 12237 4160 12287
rect 4184 12237 4219 12287
rect 4219 12237 4231 12287
rect 4231 12237 4240 12287
rect 4264 12237 4283 12287
rect 4283 12237 4320 12287
rect 3738 12231 3794 12237
rect 3818 12231 3874 12237
rect 3898 12231 3954 12237
rect 3978 12231 4034 12237
rect 4104 12231 4160 12237
rect 4184 12231 4240 12237
rect 4264 12231 4320 12237
rect 4344 12231 4400 12287
rect 3738 12147 3787 12168
rect 3787 12147 3794 12168
rect 3818 12147 3851 12168
rect 3851 12147 3863 12168
rect 3863 12147 3874 12168
rect 3898 12147 3915 12168
rect 3915 12147 3927 12168
rect 3927 12147 3954 12168
rect 3978 12147 3979 12168
rect 3979 12147 4034 12168
rect 4104 12147 4155 12168
rect 4155 12147 4160 12168
rect 4184 12147 4219 12168
rect 4219 12147 4231 12168
rect 4231 12147 4240 12168
rect 4264 12147 4283 12168
rect 4283 12147 4320 12168
rect 3738 12112 3794 12147
rect 3818 12112 3874 12147
rect 3898 12112 3954 12147
rect 3978 12112 4034 12147
rect 4104 12112 4160 12147
rect 4184 12112 4240 12147
rect 4264 12112 4320 12147
rect 4344 12112 4400 12168
rect 6468 12237 6469 12287
rect 6469 12237 6521 12287
rect 6521 12237 6524 12287
rect 6548 12237 6585 12287
rect 6585 12237 6597 12287
rect 6597 12237 6604 12287
rect 6628 12237 6649 12287
rect 6649 12237 6661 12287
rect 6661 12237 6684 12287
rect 6708 12237 6713 12287
rect 6713 12237 6764 12287
rect 6468 12231 6524 12237
rect 6548 12231 6604 12237
rect 6628 12231 6684 12237
rect 6708 12231 6764 12237
rect 6834 12237 6837 12287
rect 6837 12237 6889 12287
rect 6889 12237 6890 12287
rect 6914 12237 6953 12287
rect 6953 12237 6965 12287
rect 6965 12237 6970 12287
rect 6994 12237 7017 12287
rect 7017 12237 7050 12287
rect 6834 12231 6890 12237
rect 6914 12231 6970 12237
rect 6994 12231 7050 12237
rect 7074 12231 7130 12287
rect 6468 12147 6469 12168
rect 6469 12147 6521 12168
rect 6521 12147 6524 12168
rect 6548 12147 6585 12168
rect 6585 12147 6597 12168
rect 6597 12147 6604 12168
rect 6628 12147 6649 12168
rect 6649 12147 6661 12168
rect 6661 12147 6684 12168
rect 6708 12147 6713 12168
rect 6713 12147 6764 12168
rect 6468 12112 6524 12147
rect 6548 12112 6604 12147
rect 6628 12112 6684 12147
rect 6708 12112 6764 12147
rect 6834 12147 6837 12168
rect 6837 12147 6889 12168
rect 6889 12147 6890 12168
rect 6914 12147 6953 12168
rect 6953 12147 6965 12168
rect 6965 12147 6970 12168
rect 6994 12147 7017 12168
rect 7017 12147 7050 12168
rect 6834 12112 6890 12147
rect 6914 12112 6970 12147
rect 6994 12112 7050 12147
rect 7074 12112 7130 12168
rect 1714 12001 1770 12057
rect 1794 12001 1850 12057
rect 1874 12001 1930 12057
rect 1954 12001 2010 12057
rect 2380 12001 2436 12057
rect 2460 12001 2516 12057
rect 2540 12001 2596 12057
rect 2620 12001 2676 12057
rect 8428 12028 8484 12084
rect 8508 12028 8564 12084
rect 8588 12028 8644 12084
rect 8668 12028 8724 12084
rect 9094 12028 9150 12084
rect 9174 12028 9230 12084
rect 9254 12028 9310 12084
rect 9334 12028 9390 12084
rect 1714 11882 1770 11938
rect 1794 11882 1850 11938
rect 1874 11882 1930 11938
rect 1954 11882 2010 11938
rect 2380 11882 2436 11938
rect 2460 11882 2516 11938
rect 2540 11882 2596 11938
rect 2620 11882 2676 11938
rect 8428 11909 8484 11965
rect 8508 11909 8564 11965
rect 8588 11909 8644 11965
rect 8668 11909 8724 11965
rect 9094 11909 9150 11965
rect 9174 11909 9230 11965
rect 9254 11909 9310 11965
rect 9334 11909 9390 11965
rect 1714 181 1770 237
rect 1794 181 1850 237
rect 1874 181 1930 237
rect 1954 181 2010 237
rect 2380 181 2436 237
rect 2460 181 2516 237
rect 2540 181 2596 237
rect 2620 181 2676 237
rect 8428 188 8484 244
rect 8508 188 8564 244
rect 8588 188 8644 244
rect 8668 188 8724 244
rect 9094 188 9150 244
rect 9174 188 9230 244
rect 9254 188 9310 244
rect 9334 188 9390 244
rect 1714 62 1770 118
rect 1794 62 1850 118
rect 1874 62 1930 118
rect 1954 62 2010 118
rect 2380 62 2436 118
rect 2460 62 2516 118
rect 2540 62 2596 118
rect 2620 62 2676 118
rect 8428 69 8484 125
rect 8508 69 8564 125
rect 8588 69 8644 125
rect 8668 69 8724 125
rect 9094 69 9150 125
rect 9174 69 9230 125
rect 9254 69 9310 125
rect 9334 69 9390 125
<< metal3 >>
rect 3723 12291 4480 12296
rect 3723 12227 3734 12291
rect 3798 12227 3814 12291
rect 3878 12227 3894 12291
rect 3958 12227 3974 12291
rect 4038 12227 4100 12291
rect 4164 12227 4180 12291
rect 4244 12227 4260 12291
rect 4324 12227 4340 12291
rect 4404 12227 4480 12291
rect 1699 12061 2699 12215
rect 3723 12172 4480 12227
rect 3723 12108 3734 12172
rect 3798 12108 3814 12172
rect 3878 12108 3894 12172
rect 3958 12108 3974 12172
rect 4038 12108 4100 12172
rect 4164 12108 4180 12172
rect 4244 12108 4260 12172
rect 4324 12108 4340 12172
rect 4404 12108 4480 12172
rect 3723 12096 4480 12108
rect 6453 12291 7210 12296
rect 6453 12227 6464 12291
rect 6528 12227 6544 12291
rect 6608 12227 6624 12291
rect 6688 12227 6704 12291
rect 6768 12227 6830 12291
rect 6894 12227 6910 12291
rect 6974 12227 6990 12291
rect 7054 12227 7070 12291
rect 7134 12227 7210 12291
rect 6453 12172 7210 12227
rect 6453 12108 6464 12172
rect 6528 12108 6544 12172
rect 6608 12108 6624 12172
rect 6688 12108 6704 12172
rect 6768 12108 6830 12172
rect 6894 12108 6910 12172
rect 6974 12108 6990 12172
rect 7054 12108 7070 12172
rect 7134 12108 7210 12172
rect 6453 12096 7210 12108
rect 1699 11997 1710 12061
rect 1774 11997 1790 12061
rect 1854 11997 1870 12061
rect 1934 11997 1950 12061
rect 2014 11997 2376 12061
rect 2440 11997 2456 12061
rect 2520 11997 2536 12061
rect 2600 11997 2616 12061
rect 2680 11997 2699 12061
rect 1699 11942 2699 11997
rect 1699 11878 1710 11942
rect 1774 11878 1790 11942
rect 1854 11878 1870 11942
rect 1934 11878 1950 11942
rect 2014 11878 2376 11942
rect 2440 11878 2456 11942
rect 2520 11878 2536 11942
rect 2600 11878 2616 11942
rect 2680 11878 2699 11942
rect 8413 12088 9413 12235
rect 8413 12024 8424 12088
rect 8488 12024 8504 12088
rect 8568 12024 8584 12088
rect 8648 12024 8664 12088
rect 8728 12024 9090 12088
rect 9154 12024 9170 12088
rect 9234 12024 9250 12088
rect 9314 12024 9330 12088
rect 9394 12024 9413 12088
rect 8413 11969 9413 12024
rect 8413 11905 8424 11969
rect 8488 11905 8504 11969
rect 8568 11905 8584 11969
rect 8648 11905 8664 11969
rect 8728 11905 9090 11969
rect 9154 11905 9170 11969
rect 9234 11905 9250 11969
rect 9314 11905 9330 11969
rect 9394 11905 9413 11969
rect 8413 11893 9413 11905
rect 1699 11873 2699 11878
rect 1699 241 2699 395
rect 1699 177 1710 241
rect 1774 177 1790 241
rect 1854 177 1870 241
rect 1934 177 1950 241
rect 2014 177 2376 241
rect 2440 177 2456 241
rect 2520 177 2536 241
rect 2600 177 2616 241
rect 2680 177 2699 241
rect 1699 122 2699 177
rect 1699 58 1710 122
rect 1774 58 1790 122
rect 1854 58 1870 122
rect 1934 58 1950 122
rect 2014 58 2376 122
rect 2440 58 2456 122
rect 2520 58 2536 122
rect 2600 58 2616 122
rect 2680 58 2699 122
rect 1699 53 2699 58
rect 8413 248 9413 395
rect 8413 184 8424 248
rect 8488 184 8504 248
rect 8568 184 8584 248
rect 8648 184 8664 248
rect 8728 184 9090 248
rect 9154 184 9170 248
rect 9234 184 9250 248
rect 9314 184 9330 248
rect 9394 184 9413 248
rect 8413 129 9413 184
rect 8413 65 8424 129
rect 8488 65 8504 129
rect 8568 65 8584 129
rect 8648 65 8664 129
rect 8728 65 9090 129
rect 9154 65 9170 129
rect 9234 65 9250 129
rect 9314 65 9330 129
rect 9394 65 9413 129
rect 8413 53 9413 65
<< via3 >>
rect 3734 12287 3798 12291
rect 3734 12231 3738 12287
rect 3738 12231 3794 12287
rect 3794 12231 3798 12287
rect 3734 12227 3798 12231
rect 3814 12287 3878 12291
rect 3814 12231 3818 12287
rect 3818 12231 3874 12287
rect 3874 12231 3878 12287
rect 3814 12227 3878 12231
rect 3894 12287 3958 12291
rect 3894 12231 3898 12287
rect 3898 12231 3954 12287
rect 3954 12231 3958 12287
rect 3894 12227 3958 12231
rect 3974 12287 4038 12291
rect 3974 12231 3978 12287
rect 3978 12231 4034 12287
rect 4034 12231 4038 12287
rect 3974 12227 4038 12231
rect 4100 12287 4164 12291
rect 4100 12231 4104 12287
rect 4104 12231 4160 12287
rect 4160 12231 4164 12287
rect 4100 12227 4164 12231
rect 4180 12287 4244 12291
rect 4180 12231 4184 12287
rect 4184 12231 4240 12287
rect 4240 12231 4244 12287
rect 4180 12227 4244 12231
rect 4260 12287 4324 12291
rect 4260 12231 4264 12287
rect 4264 12231 4320 12287
rect 4320 12231 4324 12287
rect 4260 12227 4324 12231
rect 4340 12287 4404 12291
rect 4340 12231 4344 12287
rect 4344 12231 4400 12287
rect 4400 12231 4404 12287
rect 4340 12227 4404 12231
rect 3734 12168 3798 12172
rect 3734 12112 3738 12168
rect 3738 12112 3794 12168
rect 3794 12112 3798 12168
rect 3734 12108 3798 12112
rect 3814 12168 3878 12172
rect 3814 12112 3818 12168
rect 3818 12112 3874 12168
rect 3874 12112 3878 12168
rect 3814 12108 3878 12112
rect 3894 12168 3958 12172
rect 3894 12112 3898 12168
rect 3898 12112 3954 12168
rect 3954 12112 3958 12168
rect 3894 12108 3958 12112
rect 3974 12168 4038 12172
rect 3974 12112 3978 12168
rect 3978 12112 4034 12168
rect 4034 12112 4038 12168
rect 3974 12108 4038 12112
rect 4100 12168 4164 12172
rect 4100 12112 4104 12168
rect 4104 12112 4160 12168
rect 4160 12112 4164 12168
rect 4100 12108 4164 12112
rect 4180 12168 4244 12172
rect 4180 12112 4184 12168
rect 4184 12112 4240 12168
rect 4240 12112 4244 12168
rect 4180 12108 4244 12112
rect 4260 12168 4324 12172
rect 4260 12112 4264 12168
rect 4264 12112 4320 12168
rect 4320 12112 4324 12168
rect 4260 12108 4324 12112
rect 4340 12168 4404 12172
rect 4340 12112 4344 12168
rect 4344 12112 4400 12168
rect 4400 12112 4404 12168
rect 4340 12108 4404 12112
rect 6464 12287 6528 12291
rect 6464 12231 6468 12287
rect 6468 12231 6524 12287
rect 6524 12231 6528 12287
rect 6464 12227 6528 12231
rect 6544 12287 6608 12291
rect 6544 12231 6548 12287
rect 6548 12231 6604 12287
rect 6604 12231 6608 12287
rect 6544 12227 6608 12231
rect 6624 12287 6688 12291
rect 6624 12231 6628 12287
rect 6628 12231 6684 12287
rect 6684 12231 6688 12287
rect 6624 12227 6688 12231
rect 6704 12287 6768 12291
rect 6704 12231 6708 12287
rect 6708 12231 6764 12287
rect 6764 12231 6768 12287
rect 6704 12227 6768 12231
rect 6830 12287 6894 12291
rect 6830 12231 6834 12287
rect 6834 12231 6890 12287
rect 6890 12231 6894 12287
rect 6830 12227 6894 12231
rect 6910 12287 6974 12291
rect 6910 12231 6914 12287
rect 6914 12231 6970 12287
rect 6970 12231 6974 12287
rect 6910 12227 6974 12231
rect 6990 12287 7054 12291
rect 6990 12231 6994 12287
rect 6994 12231 7050 12287
rect 7050 12231 7054 12287
rect 6990 12227 7054 12231
rect 7070 12287 7134 12291
rect 7070 12231 7074 12287
rect 7074 12231 7130 12287
rect 7130 12231 7134 12287
rect 7070 12227 7134 12231
rect 6464 12168 6528 12172
rect 6464 12112 6468 12168
rect 6468 12112 6524 12168
rect 6524 12112 6528 12168
rect 6464 12108 6528 12112
rect 6544 12168 6608 12172
rect 6544 12112 6548 12168
rect 6548 12112 6604 12168
rect 6604 12112 6608 12168
rect 6544 12108 6608 12112
rect 6624 12168 6688 12172
rect 6624 12112 6628 12168
rect 6628 12112 6684 12168
rect 6684 12112 6688 12168
rect 6624 12108 6688 12112
rect 6704 12168 6768 12172
rect 6704 12112 6708 12168
rect 6708 12112 6764 12168
rect 6764 12112 6768 12168
rect 6704 12108 6768 12112
rect 6830 12168 6894 12172
rect 6830 12112 6834 12168
rect 6834 12112 6890 12168
rect 6890 12112 6894 12168
rect 6830 12108 6894 12112
rect 6910 12168 6974 12172
rect 6910 12112 6914 12168
rect 6914 12112 6970 12168
rect 6970 12112 6974 12168
rect 6910 12108 6974 12112
rect 6990 12168 7054 12172
rect 6990 12112 6994 12168
rect 6994 12112 7050 12168
rect 7050 12112 7054 12168
rect 6990 12108 7054 12112
rect 7070 12168 7134 12172
rect 7070 12112 7074 12168
rect 7074 12112 7130 12168
rect 7130 12112 7134 12168
rect 7070 12108 7134 12112
rect 1710 12057 1774 12061
rect 1710 12001 1714 12057
rect 1714 12001 1770 12057
rect 1770 12001 1774 12057
rect 1710 11997 1774 12001
rect 1790 12057 1854 12061
rect 1790 12001 1794 12057
rect 1794 12001 1850 12057
rect 1850 12001 1854 12057
rect 1790 11997 1854 12001
rect 1870 12057 1934 12061
rect 1870 12001 1874 12057
rect 1874 12001 1930 12057
rect 1930 12001 1934 12057
rect 1870 11997 1934 12001
rect 1950 12057 2014 12061
rect 1950 12001 1954 12057
rect 1954 12001 2010 12057
rect 2010 12001 2014 12057
rect 1950 11997 2014 12001
rect 2376 12057 2440 12061
rect 2376 12001 2380 12057
rect 2380 12001 2436 12057
rect 2436 12001 2440 12057
rect 2376 11997 2440 12001
rect 2456 12057 2520 12061
rect 2456 12001 2460 12057
rect 2460 12001 2516 12057
rect 2516 12001 2520 12057
rect 2456 11997 2520 12001
rect 2536 12057 2600 12061
rect 2536 12001 2540 12057
rect 2540 12001 2596 12057
rect 2596 12001 2600 12057
rect 2536 11997 2600 12001
rect 2616 12057 2680 12061
rect 2616 12001 2620 12057
rect 2620 12001 2676 12057
rect 2676 12001 2680 12057
rect 2616 11997 2680 12001
rect 1710 11938 1774 11942
rect 1710 11882 1714 11938
rect 1714 11882 1770 11938
rect 1770 11882 1774 11938
rect 1710 11878 1774 11882
rect 1790 11938 1854 11942
rect 1790 11882 1794 11938
rect 1794 11882 1850 11938
rect 1850 11882 1854 11938
rect 1790 11878 1854 11882
rect 1870 11938 1934 11942
rect 1870 11882 1874 11938
rect 1874 11882 1930 11938
rect 1930 11882 1934 11938
rect 1870 11878 1934 11882
rect 1950 11938 2014 11942
rect 1950 11882 1954 11938
rect 1954 11882 2010 11938
rect 2010 11882 2014 11938
rect 1950 11878 2014 11882
rect 2376 11938 2440 11942
rect 2376 11882 2380 11938
rect 2380 11882 2436 11938
rect 2436 11882 2440 11938
rect 2376 11878 2440 11882
rect 2456 11938 2520 11942
rect 2456 11882 2460 11938
rect 2460 11882 2516 11938
rect 2516 11882 2520 11938
rect 2456 11878 2520 11882
rect 2536 11938 2600 11942
rect 2536 11882 2540 11938
rect 2540 11882 2596 11938
rect 2596 11882 2600 11938
rect 2536 11878 2600 11882
rect 2616 11938 2680 11942
rect 2616 11882 2620 11938
rect 2620 11882 2676 11938
rect 2676 11882 2680 11938
rect 2616 11878 2680 11882
rect 8424 12084 8488 12088
rect 8424 12028 8428 12084
rect 8428 12028 8484 12084
rect 8484 12028 8488 12084
rect 8424 12024 8488 12028
rect 8504 12084 8568 12088
rect 8504 12028 8508 12084
rect 8508 12028 8564 12084
rect 8564 12028 8568 12084
rect 8504 12024 8568 12028
rect 8584 12084 8648 12088
rect 8584 12028 8588 12084
rect 8588 12028 8644 12084
rect 8644 12028 8648 12084
rect 8584 12024 8648 12028
rect 8664 12084 8728 12088
rect 8664 12028 8668 12084
rect 8668 12028 8724 12084
rect 8724 12028 8728 12084
rect 8664 12024 8728 12028
rect 9090 12084 9154 12088
rect 9090 12028 9094 12084
rect 9094 12028 9150 12084
rect 9150 12028 9154 12084
rect 9090 12024 9154 12028
rect 9170 12084 9234 12088
rect 9170 12028 9174 12084
rect 9174 12028 9230 12084
rect 9230 12028 9234 12084
rect 9170 12024 9234 12028
rect 9250 12084 9314 12088
rect 9250 12028 9254 12084
rect 9254 12028 9310 12084
rect 9310 12028 9314 12084
rect 9250 12024 9314 12028
rect 9330 12084 9394 12088
rect 9330 12028 9334 12084
rect 9334 12028 9390 12084
rect 9390 12028 9394 12084
rect 9330 12024 9394 12028
rect 8424 11965 8488 11969
rect 8424 11909 8428 11965
rect 8428 11909 8484 11965
rect 8484 11909 8488 11965
rect 8424 11905 8488 11909
rect 8504 11965 8568 11969
rect 8504 11909 8508 11965
rect 8508 11909 8564 11965
rect 8564 11909 8568 11965
rect 8504 11905 8568 11909
rect 8584 11965 8648 11969
rect 8584 11909 8588 11965
rect 8588 11909 8644 11965
rect 8644 11909 8648 11965
rect 8584 11905 8648 11909
rect 8664 11965 8728 11969
rect 8664 11909 8668 11965
rect 8668 11909 8724 11965
rect 8724 11909 8728 11965
rect 8664 11905 8728 11909
rect 9090 11965 9154 11969
rect 9090 11909 9094 11965
rect 9094 11909 9150 11965
rect 9150 11909 9154 11965
rect 9090 11905 9154 11909
rect 9170 11965 9234 11969
rect 9170 11909 9174 11965
rect 9174 11909 9230 11965
rect 9230 11909 9234 11965
rect 9170 11905 9234 11909
rect 9250 11965 9314 11969
rect 9250 11909 9254 11965
rect 9254 11909 9310 11965
rect 9310 11909 9314 11965
rect 9250 11905 9314 11909
rect 9330 11965 9394 11969
rect 9330 11909 9334 11965
rect 9334 11909 9390 11965
rect 9390 11909 9394 11965
rect 9330 11905 9394 11909
rect 1710 237 1774 241
rect 1710 181 1714 237
rect 1714 181 1770 237
rect 1770 181 1774 237
rect 1710 177 1774 181
rect 1790 237 1854 241
rect 1790 181 1794 237
rect 1794 181 1850 237
rect 1850 181 1854 237
rect 1790 177 1854 181
rect 1870 237 1934 241
rect 1870 181 1874 237
rect 1874 181 1930 237
rect 1930 181 1934 237
rect 1870 177 1934 181
rect 1950 237 2014 241
rect 1950 181 1954 237
rect 1954 181 2010 237
rect 2010 181 2014 237
rect 1950 177 2014 181
rect 2376 237 2440 241
rect 2376 181 2380 237
rect 2380 181 2436 237
rect 2436 181 2440 237
rect 2376 177 2440 181
rect 2456 237 2520 241
rect 2456 181 2460 237
rect 2460 181 2516 237
rect 2516 181 2520 237
rect 2456 177 2520 181
rect 2536 237 2600 241
rect 2536 181 2540 237
rect 2540 181 2596 237
rect 2596 181 2600 237
rect 2536 177 2600 181
rect 2616 237 2680 241
rect 2616 181 2620 237
rect 2620 181 2676 237
rect 2676 181 2680 237
rect 2616 177 2680 181
rect 1710 118 1774 122
rect 1710 62 1714 118
rect 1714 62 1770 118
rect 1770 62 1774 118
rect 1710 58 1774 62
rect 1790 118 1854 122
rect 1790 62 1794 118
rect 1794 62 1850 118
rect 1850 62 1854 118
rect 1790 58 1854 62
rect 1870 118 1934 122
rect 1870 62 1874 118
rect 1874 62 1930 118
rect 1930 62 1934 118
rect 1870 58 1934 62
rect 1950 118 2014 122
rect 1950 62 1954 118
rect 1954 62 2010 118
rect 2010 62 2014 118
rect 1950 58 2014 62
rect 2376 118 2440 122
rect 2376 62 2380 118
rect 2380 62 2436 118
rect 2436 62 2440 118
rect 2376 58 2440 62
rect 2456 118 2520 122
rect 2456 62 2460 118
rect 2460 62 2516 118
rect 2516 62 2520 118
rect 2456 58 2520 62
rect 2536 118 2600 122
rect 2536 62 2540 118
rect 2540 62 2596 118
rect 2596 62 2600 118
rect 2536 58 2600 62
rect 2616 118 2680 122
rect 2616 62 2620 118
rect 2620 62 2676 118
rect 2676 62 2680 118
rect 2616 58 2680 62
rect 8424 244 8488 248
rect 8424 188 8428 244
rect 8428 188 8484 244
rect 8484 188 8488 244
rect 8424 184 8488 188
rect 8504 244 8568 248
rect 8504 188 8508 244
rect 8508 188 8564 244
rect 8564 188 8568 244
rect 8504 184 8568 188
rect 8584 244 8648 248
rect 8584 188 8588 244
rect 8588 188 8644 244
rect 8644 188 8648 244
rect 8584 184 8648 188
rect 8664 244 8728 248
rect 8664 188 8668 244
rect 8668 188 8724 244
rect 8724 188 8728 244
rect 8664 184 8728 188
rect 9090 244 9154 248
rect 9090 188 9094 244
rect 9094 188 9150 244
rect 9150 188 9154 244
rect 9090 184 9154 188
rect 9170 244 9234 248
rect 9170 188 9174 244
rect 9174 188 9230 244
rect 9230 188 9234 244
rect 9170 184 9234 188
rect 9250 244 9314 248
rect 9250 188 9254 244
rect 9254 188 9310 244
rect 9310 188 9314 244
rect 9250 184 9314 188
rect 9330 244 9394 248
rect 9330 188 9334 244
rect 9334 188 9390 244
rect 9390 188 9394 244
rect 9330 184 9394 188
rect 8424 125 8488 129
rect 8424 69 8428 125
rect 8428 69 8484 125
rect 8484 69 8488 125
rect 8424 65 8488 69
rect 8504 125 8568 129
rect 8504 69 8508 125
rect 8508 69 8564 125
rect 8564 69 8568 125
rect 8504 65 8568 69
rect 8584 125 8648 129
rect 8584 69 8588 125
rect 8588 69 8644 125
rect 8644 69 8648 125
rect 8584 65 8648 69
rect 8664 125 8728 129
rect 8664 69 8668 125
rect 8668 69 8724 125
rect 8724 69 8728 125
rect 8664 65 8728 69
rect 9090 125 9154 129
rect 9090 69 9094 125
rect 9094 69 9150 125
rect 9150 69 9154 125
rect 9090 65 9154 69
rect 9170 125 9234 129
rect 9170 69 9174 125
rect 9174 69 9230 125
rect 9230 69 9234 125
rect 9170 65 9234 69
rect 9250 125 9314 129
rect 9250 69 9254 125
rect 9254 69 9310 125
rect 9310 69 9314 125
rect 9250 65 9314 69
rect 9330 125 9394 129
rect 9330 69 9334 125
rect 9334 69 9390 125
rect 9390 69 9394 125
rect 9330 65 9394 69
<< metal4 >>
rect 1699 12061 2699 18646
rect 3723 12291 4480 19729
rect 3723 12227 3734 12291
rect 3798 12227 3814 12291
rect 3878 12227 3894 12291
rect 3958 12227 3974 12291
rect 4038 12227 4100 12291
rect 4164 12227 4180 12291
rect 4244 12227 4260 12291
rect 4324 12227 4340 12291
rect 4404 12227 4480 12291
rect 3723 12172 4480 12227
rect 3723 12108 3734 12172
rect 3798 12108 3814 12172
rect 3878 12108 3894 12172
rect 3958 12108 3974 12172
rect 4038 12108 4100 12172
rect 4164 12108 4180 12172
rect 4244 12108 4260 12172
rect 4324 12108 4340 12172
rect 4404 12108 4480 12172
rect 3723 12096 4480 12108
rect 6453 12291 7210 19729
rect 6453 12227 6464 12291
rect 6528 12227 6544 12291
rect 6608 12227 6624 12291
rect 6688 12227 6704 12291
rect 6768 12227 6830 12291
rect 6894 12227 6910 12291
rect 6974 12227 6990 12291
rect 7054 12227 7070 12291
rect 7134 12227 7210 12291
rect 6453 12172 7210 12227
rect 6453 12108 6464 12172
rect 6528 12108 6544 12172
rect 6608 12108 6624 12172
rect 6688 12108 6704 12172
rect 6768 12108 6830 12172
rect 6894 12108 6910 12172
rect 6974 12108 6990 12172
rect 7054 12108 7070 12172
rect 7134 12108 7210 12172
rect 6453 12096 7210 12108
rect 1699 11997 1710 12061
rect 1774 11997 1790 12061
rect 1854 11997 1870 12061
rect 1934 11997 1950 12061
rect 2014 11997 2376 12061
rect 2440 11997 2456 12061
rect 2520 11997 2536 12061
rect 2600 11997 2616 12061
rect 2680 11997 2699 12061
rect 1699 11942 2699 11997
rect 1699 11878 1710 11942
rect 1774 11878 1790 11942
rect 1854 11878 1870 11942
rect 1934 11878 1950 11942
rect 2014 11878 2376 11942
rect 2440 11878 2456 11942
rect 2520 11878 2536 11942
rect 2600 11878 2616 11942
rect 2680 11878 2699 11942
rect 1699 241 2699 11878
rect 1699 177 1710 241
rect 1774 177 1790 241
rect 1854 177 1870 241
rect 1934 177 1950 241
rect 2014 177 2376 241
rect 2440 177 2456 241
rect 2520 177 2536 241
rect 2600 177 2616 241
rect 2680 177 2699 241
rect 1699 122 2699 177
rect 1699 58 1710 122
rect 1774 58 1790 122
rect 1854 58 1870 122
rect 1934 58 1950 122
rect 2014 58 2376 122
rect 2440 58 2456 122
rect 2520 58 2536 122
rect 2600 58 2616 122
rect 2680 58 2699 122
rect 1699 -6410 2699 58
rect 8413 12088 9413 18646
rect 8413 12024 8424 12088
rect 8488 12024 8504 12088
rect 8568 12024 8584 12088
rect 8648 12024 8664 12088
rect 8728 12024 9090 12088
rect 9154 12024 9170 12088
rect 9234 12024 9250 12088
rect 9314 12024 9330 12088
rect 9394 12024 9413 12088
rect 8413 11969 9413 12024
rect 8413 11905 8424 11969
rect 8488 11905 8504 11969
rect 8568 11905 8584 11969
rect 8648 11905 8664 11969
rect 8728 11905 9090 11969
rect 9154 11905 9170 11969
rect 9234 11905 9250 11969
rect 9314 11905 9330 11969
rect 9394 11905 9413 11969
rect 8413 248 9413 11905
rect 8413 184 8424 248
rect 8488 184 8504 248
rect 8568 184 8584 248
rect 8648 184 8664 248
rect 8728 184 9090 248
rect 9154 184 9170 248
rect 9234 184 9250 248
rect 9314 184 9330 248
rect 9394 184 9413 248
rect 8413 129 9413 184
rect 8413 65 8424 129
rect 8488 65 8504 129
rect 8568 65 8584 129
rect 8648 65 8664 129
rect 8728 65 9090 129
rect 9154 65 9170 129
rect 9234 65 9250 129
rect 9314 65 9330 129
rect 9394 65 9413 129
rect 8413 -6410 9413 65
use sky130_ef_ip__rc_osc_500k  sky130_ef_ip__rc_osc_500k_0
timestamp 1528465711
transform 0 -1 10844 1 0 54
box 0 0 12242 10724
<< labels >>
flabel metal2 s 5933 12473 6045 13913 0 FreeSans 560 90 0 0 ena
port 1 nsew
flabel metal2 s 5289 12473 5401 13913 0 FreeSans 560 90 0 0 dout
port 2 nsew
flabel metal4 s 8413 -6410 9413 18646 0 FreeSans 9600 90 0 0 vssa1
port 3 nsew
flabel metal4 s 1699 -6410 2699 18646 0 FreeSans 9600 90 0 0 vdda1
port 4 nsew
flabel metal4 s 6453 12096 7210 19729 0 FreeSans 9600 90 0 0 vccd1
port 5 nsew
flabel metal4 s 3723 12096 4480 19729 0 FreeSans 9600 90 0 0 vssd1
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 10872 12778
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1527881472
<< checkpaint >>
rect -4796 -3724 23196 23852
<< metal2 >>
rect 9006 20210 9118 21516
rect 9650 20316 9762 21516
rect 8864 20182 9118 20210
rect 7440 16233 8197 16242
rect 7440 16177 7455 16233
rect 7511 16177 7535 16233
rect 7591 16177 7615 16233
rect 7671 16177 7695 16233
rect 7751 16177 7821 16233
rect 7877 16177 7901 16233
rect 7957 16177 7981 16233
rect 8037 16177 8061 16233
rect 8117 16177 8197 16233
rect 7440 16114 8197 16177
rect 8864 16116 8892 20182
rect 9006 20076 9118 20182
rect 9641 20076 9762 20316
rect 9641 20074 9669 20076
rect 9600 20046 9669 20074
rect 9600 16116 9628 20046
rect 10170 16233 10927 16242
rect 10170 16177 10185 16233
rect 10241 16177 10265 16233
rect 10321 16177 10345 16233
rect 10401 16177 10425 16233
rect 10481 16177 10551 16233
rect 10607 16177 10631 16233
rect 10687 16177 10711 16233
rect 10767 16177 10791 16233
rect 10847 16177 10927 16233
rect 7440 16058 7455 16114
rect 7511 16058 7535 16114
rect 7591 16058 7615 16114
rect 7671 16058 7695 16114
rect 7751 16058 7821 16114
rect 7877 16058 7901 16114
rect 7957 16058 7981 16114
rect 8037 16058 8061 16114
rect 8117 16058 8197 16114
rect 7440 16042 8197 16058
rect 10170 16114 10927 16177
rect 10170 16058 10185 16114
rect 10241 16058 10265 16114
rect 10321 16058 10345 16114
rect 10401 16058 10425 16114
rect 10481 16058 10551 16114
rect 10607 16058 10631 16114
rect 10687 16058 10711 16114
rect 10767 16058 10791 16114
rect 10847 16058 10927 16114
rect 10170 16042 10927 16058
<< via2 >>
rect 7455 16177 7511 16233
rect 7535 16177 7591 16233
rect 7615 16177 7671 16233
rect 7695 16177 7751 16233
rect 7821 16177 7877 16233
rect 7901 16177 7957 16233
rect 7981 16177 8037 16233
rect 8061 16177 8117 16233
rect 10185 16177 10241 16233
rect 10265 16177 10321 16233
rect 10345 16177 10401 16233
rect 10425 16177 10481 16233
rect 10551 16177 10607 16233
rect 10631 16177 10687 16233
rect 10711 16177 10767 16233
rect 10791 16177 10847 16233
rect 7455 16058 7511 16114
rect 7535 16058 7591 16114
rect 7615 16058 7671 16114
rect 7695 16058 7751 16114
rect 7821 16058 7877 16114
rect 7901 16058 7957 16114
rect 7981 16058 8037 16114
rect 8061 16058 8117 16114
rect 10185 16058 10241 16114
rect 10265 16058 10321 16114
rect 10345 16058 10401 16114
rect 10425 16058 10481 16114
rect 10551 16058 10607 16114
rect 10631 16058 10687 16114
rect 10711 16058 10767 16114
rect 10791 16058 10847 16114
rect 5431 4127 5487 4183
rect 5511 4127 5567 4183
rect 5591 4127 5647 4183
rect 5671 4127 5727 4183
rect 6097 4127 6153 4183
rect 6177 4127 6233 4183
rect 6257 4127 6313 4183
rect 6337 4127 6393 4183
rect 12145 4134 12201 4190
rect 12225 4134 12281 4190
rect 12305 4134 12361 4190
rect 12385 4134 12441 4190
rect 12811 4134 12867 4190
rect 12891 4134 12947 4190
rect 12971 4134 13027 4190
rect 13051 4134 13107 4190
rect 5431 4008 5487 4064
rect 5511 4008 5567 4064
rect 5591 4008 5647 4064
rect 5671 4008 5727 4064
rect 6097 4008 6153 4064
rect 6177 4008 6233 4064
rect 6257 4008 6313 4064
rect 6337 4008 6393 4064
rect 12145 4015 12201 4071
rect 12225 4015 12281 4071
rect 12305 4015 12361 4071
rect 12385 4015 12441 4071
rect 12811 4015 12867 4071
rect 12891 4015 12947 4071
rect 12971 4015 13027 4071
rect 13051 4015 13107 4071
<< metal3 >>
rect 7440 16237 8197 16242
rect 7440 16173 7451 16237
rect 7515 16173 7531 16237
rect 7595 16173 7611 16237
rect 7675 16173 7691 16237
rect 7755 16173 7817 16237
rect 7881 16173 7897 16237
rect 7961 16173 7977 16237
rect 8041 16173 8057 16237
rect 8121 16173 8197 16237
rect 7440 16118 8197 16173
rect 7440 16054 7451 16118
rect 7515 16054 7531 16118
rect 7595 16054 7611 16118
rect 7675 16054 7691 16118
rect 7755 16054 7817 16118
rect 7881 16054 7897 16118
rect 7961 16054 7977 16118
rect 8041 16054 8057 16118
rect 8121 16054 8197 16118
rect 7440 16042 8197 16054
rect 10170 16237 10927 16242
rect 10170 16173 10181 16237
rect 10245 16173 10261 16237
rect 10325 16173 10341 16237
rect 10405 16173 10421 16237
rect 10485 16173 10547 16237
rect 10611 16173 10627 16237
rect 10691 16173 10707 16237
rect 10771 16173 10787 16237
rect 10851 16173 10927 16237
rect 10170 16118 10927 16173
rect 10170 16054 10181 16118
rect 10245 16054 10261 16118
rect 10325 16054 10341 16118
rect 10405 16054 10421 16118
rect 10485 16054 10547 16118
rect 10611 16054 10627 16118
rect 10691 16054 10707 16118
rect 10771 16054 10787 16118
rect 10851 16054 10927 16118
rect 10170 16042 10927 16054
rect 5416 4187 6416 4341
rect 5416 4123 5427 4187
rect 5491 4123 5507 4187
rect 5571 4123 5587 4187
rect 5651 4123 5667 4187
rect 5731 4123 6093 4187
rect 6157 4123 6173 4187
rect 6237 4123 6253 4187
rect 6317 4123 6333 4187
rect 6397 4123 6416 4187
rect 5416 4068 6416 4123
rect 5416 4004 5427 4068
rect 5491 4004 5507 4068
rect 5571 4004 5587 4068
rect 5651 4004 5667 4068
rect 5731 4004 6093 4068
rect 6157 4004 6173 4068
rect 6237 4004 6253 4068
rect 6317 4004 6333 4068
rect 6397 4004 6416 4068
rect 5416 3999 6416 4004
rect 12130 4194 13130 4341
rect 12130 4130 12141 4194
rect 12205 4130 12221 4194
rect 12285 4130 12301 4194
rect 12365 4130 12381 4194
rect 12445 4130 12807 4194
rect 12871 4130 12887 4194
rect 12951 4130 12967 4194
rect 13031 4130 13047 4194
rect 13111 4130 13130 4194
rect 12130 4075 13130 4130
rect 12130 4011 12141 4075
rect 12205 4011 12221 4075
rect 12285 4011 12301 4075
rect 12365 4011 12381 4075
rect 12445 4011 12807 4075
rect 12871 4011 12887 4075
rect 12951 4011 12967 4075
rect 13031 4011 13047 4075
rect 13111 4011 13130 4075
rect 12130 3999 13130 4011
<< via3 >>
rect 7451 16233 7515 16237
rect 7451 16177 7455 16233
rect 7455 16177 7511 16233
rect 7511 16177 7515 16233
rect 7451 16173 7515 16177
rect 7531 16233 7595 16237
rect 7531 16177 7535 16233
rect 7535 16177 7591 16233
rect 7591 16177 7595 16233
rect 7531 16173 7595 16177
rect 7611 16233 7675 16237
rect 7611 16177 7615 16233
rect 7615 16177 7671 16233
rect 7671 16177 7675 16233
rect 7611 16173 7675 16177
rect 7691 16233 7755 16237
rect 7691 16177 7695 16233
rect 7695 16177 7751 16233
rect 7751 16177 7755 16233
rect 7691 16173 7755 16177
rect 7817 16233 7881 16237
rect 7817 16177 7821 16233
rect 7821 16177 7877 16233
rect 7877 16177 7881 16233
rect 7817 16173 7881 16177
rect 7897 16233 7961 16237
rect 7897 16177 7901 16233
rect 7901 16177 7957 16233
rect 7957 16177 7961 16233
rect 7897 16173 7961 16177
rect 7977 16233 8041 16237
rect 7977 16177 7981 16233
rect 7981 16177 8037 16233
rect 8037 16177 8041 16233
rect 7977 16173 8041 16177
rect 8057 16233 8121 16237
rect 8057 16177 8061 16233
rect 8061 16177 8117 16233
rect 8117 16177 8121 16233
rect 8057 16173 8121 16177
rect 7451 16114 7515 16118
rect 7451 16058 7455 16114
rect 7455 16058 7511 16114
rect 7511 16058 7515 16114
rect 7451 16054 7515 16058
rect 7531 16114 7595 16118
rect 7531 16058 7535 16114
rect 7535 16058 7591 16114
rect 7591 16058 7595 16114
rect 7531 16054 7595 16058
rect 7611 16114 7675 16118
rect 7611 16058 7615 16114
rect 7615 16058 7671 16114
rect 7671 16058 7675 16114
rect 7611 16054 7675 16058
rect 7691 16114 7755 16118
rect 7691 16058 7695 16114
rect 7695 16058 7751 16114
rect 7751 16058 7755 16114
rect 7691 16054 7755 16058
rect 7817 16114 7881 16118
rect 7817 16058 7821 16114
rect 7821 16058 7877 16114
rect 7877 16058 7881 16114
rect 7817 16054 7881 16058
rect 7897 16114 7961 16118
rect 7897 16058 7901 16114
rect 7901 16058 7957 16114
rect 7957 16058 7961 16114
rect 7897 16054 7961 16058
rect 7977 16114 8041 16118
rect 7977 16058 7981 16114
rect 7981 16058 8037 16114
rect 8037 16058 8041 16114
rect 7977 16054 8041 16058
rect 8057 16114 8121 16118
rect 8057 16058 8061 16114
rect 8061 16058 8117 16114
rect 8117 16058 8121 16114
rect 8057 16054 8121 16058
rect 10181 16233 10245 16237
rect 10181 16177 10185 16233
rect 10185 16177 10241 16233
rect 10241 16177 10245 16233
rect 10181 16173 10245 16177
rect 10261 16233 10325 16237
rect 10261 16177 10265 16233
rect 10265 16177 10321 16233
rect 10321 16177 10325 16233
rect 10261 16173 10325 16177
rect 10341 16233 10405 16237
rect 10341 16177 10345 16233
rect 10345 16177 10401 16233
rect 10401 16177 10405 16233
rect 10341 16173 10405 16177
rect 10421 16233 10485 16237
rect 10421 16177 10425 16233
rect 10425 16177 10481 16233
rect 10481 16177 10485 16233
rect 10421 16173 10485 16177
rect 10547 16233 10611 16237
rect 10547 16177 10551 16233
rect 10551 16177 10607 16233
rect 10607 16177 10611 16233
rect 10547 16173 10611 16177
rect 10627 16233 10691 16237
rect 10627 16177 10631 16233
rect 10631 16177 10687 16233
rect 10687 16177 10691 16233
rect 10627 16173 10691 16177
rect 10707 16233 10771 16237
rect 10707 16177 10711 16233
rect 10711 16177 10767 16233
rect 10767 16177 10771 16233
rect 10707 16173 10771 16177
rect 10787 16233 10851 16237
rect 10787 16177 10791 16233
rect 10791 16177 10847 16233
rect 10847 16177 10851 16233
rect 10787 16173 10851 16177
rect 10181 16114 10245 16118
rect 10181 16058 10185 16114
rect 10185 16058 10241 16114
rect 10241 16058 10245 16114
rect 10181 16054 10245 16058
rect 10261 16114 10325 16118
rect 10261 16058 10265 16114
rect 10265 16058 10321 16114
rect 10321 16058 10325 16114
rect 10261 16054 10325 16058
rect 10341 16114 10405 16118
rect 10341 16058 10345 16114
rect 10345 16058 10401 16114
rect 10401 16058 10405 16114
rect 10341 16054 10405 16058
rect 10421 16114 10485 16118
rect 10421 16058 10425 16114
rect 10425 16058 10481 16114
rect 10481 16058 10485 16114
rect 10421 16054 10485 16058
rect 10547 16114 10611 16118
rect 10547 16058 10551 16114
rect 10551 16058 10607 16114
rect 10607 16058 10611 16114
rect 10547 16054 10611 16058
rect 10627 16114 10691 16118
rect 10627 16058 10631 16114
rect 10631 16058 10687 16114
rect 10687 16058 10691 16114
rect 10627 16054 10691 16058
rect 10707 16114 10771 16118
rect 10707 16058 10711 16114
rect 10711 16058 10767 16114
rect 10767 16058 10771 16114
rect 10707 16054 10771 16058
rect 10787 16114 10851 16118
rect 10787 16058 10791 16114
rect 10791 16058 10847 16114
rect 10847 16058 10851 16114
rect 10787 16054 10851 16058
rect 5427 4183 5491 4187
rect 5427 4127 5431 4183
rect 5431 4127 5487 4183
rect 5487 4127 5491 4183
rect 5427 4123 5491 4127
rect 5507 4183 5571 4187
rect 5507 4127 5511 4183
rect 5511 4127 5567 4183
rect 5567 4127 5571 4183
rect 5507 4123 5571 4127
rect 5587 4183 5651 4187
rect 5587 4127 5591 4183
rect 5591 4127 5647 4183
rect 5647 4127 5651 4183
rect 5587 4123 5651 4127
rect 5667 4183 5731 4187
rect 5667 4127 5671 4183
rect 5671 4127 5727 4183
rect 5727 4127 5731 4183
rect 5667 4123 5731 4127
rect 6093 4183 6157 4187
rect 6093 4127 6097 4183
rect 6097 4127 6153 4183
rect 6153 4127 6157 4183
rect 6093 4123 6157 4127
rect 6173 4183 6237 4187
rect 6173 4127 6177 4183
rect 6177 4127 6233 4183
rect 6233 4127 6237 4183
rect 6173 4123 6237 4127
rect 6253 4183 6317 4187
rect 6253 4127 6257 4183
rect 6257 4127 6313 4183
rect 6313 4127 6317 4183
rect 6253 4123 6317 4127
rect 6333 4183 6397 4187
rect 6333 4127 6337 4183
rect 6337 4127 6393 4183
rect 6393 4127 6397 4183
rect 6333 4123 6397 4127
rect 5427 4064 5491 4068
rect 5427 4008 5431 4064
rect 5431 4008 5487 4064
rect 5487 4008 5491 4064
rect 5427 4004 5491 4008
rect 5507 4064 5571 4068
rect 5507 4008 5511 4064
rect 5511 4008 5567 4064
rect 5567 4008 5571 4064
rect 5507 4004 5571 4008
rect 5587 4064 5651 4068
rect 5587 4008 5591 4064
rect 5591 4008 5647 4064
rect 5647 4008 5651 4064
rect 5587 4004 5651 4008
rect 5667 4064 5731 4068
rect 5667 4008 5671 4064
rect 5671 4008 5727 4064
rect 5727 4008 5731 4064
rect 5667 4004 5731 4008
rect 6093 4064 6157 4068
rect 6093 4008 6097 4064
rect 6097 4008 6153 4064
rect 6153 4008 6157 4064
rect 6093 4004 6157 4008
rect 6173 4064 6237 4068
rect 6173 4008 6177 4064
rect 6177 4008 6233 4064
rect 6233 4008 6237 4064
rect 6173 4004 6237 4008
rect 6253 4064 6317 4068
rect 6253 4008 6257 4064
rect 6257 4008 6313 4064
rect 6313 4008 6317 4064
rect 6253 4004 6317 4008
rect 6333 4064 6397 4068
rect 6333 4008 6337 4064
rect 6337 4008 6393 4064
rect 6393 4008 6397 4064
rect 6333 4004 6397 4008
rect 12141 4190 12205 4194
rect 12141 4134 12145 4190
rect 12145 4134 12201 4190
rect 12201 4134 12205 4190
rect 12141 4130 12205 4134
rect 12221 4190 12285 4194
rect 12221 4134 12225 4190
rect 12225 4134 12281 4190
rect 12281 4134 12285 4190
rect 12221 4130 12285 4134
rect 12301 4190 12365 4194
rect 12301 4134 12305 4190
rect 12305 4134 12361 4190
rect 12361 4134 12365 4190
rect 12301 4130 12365 4134
rect 12381 4190 12445 4194
rect 12381 4134 12385 4190
rect 12385 4134 12441 4190
rect 12441 4134 12445 4190
rect 12381 4130 12445 4134
rect 12807 4190 12871 4194
rect 12807 4134 12811 4190
rect 12811 4134 12867 4190
rect 12867 4134 12871 4190
rect 12807 4130 12871 4134
rect 12887 4190 12951 4194
rect 12887 4134 12891 4190
rect 12891 4134 12947 4190
rect 12947 4134 12951 4190
rect 12887 4130 12951 4134
rect 12967 4190 13031 4194
rect 12967 4134 12971 4190
rect 12971 4134 13027 4190
rect 13027 4134 13031 4190
rect 12967 4130 13031 4134
rect 13047 4190 13111 4194
rect 13047 4134 13051 4190
rect 13051 4134 13107 4190
rect 13107 4134 13111 4190
rect 13047 4130 13111 4134
rect 12141 4071 12205 4075
rect 12141 4015 12145 4071
rect 12145 4015 12201 4071
rect 12201 4015 12205 4071
rect 12141 4011 12205 4015
rect 12221 4071 12285 4075
rect 12221 4015 12225 4071
rect 12225 4015 12281 4071
rect 12281 4015 12285 4071
rect 12221 4011 12285 4015
rect 12301 4071 12365 4075
rect 12301 4015 12305 4071
rect 12305 4015 12361 4071
rect 12361 4015 12365 4071
rect 12301 4011 12365 4015
rect 12381 4071 12445 4075
rect 12381 4015 12385 4071
rect 12385 4015 12441 4071
rect 12441 4015 12445 4071
rect 12381 4011 12445 4015
rect 12807 4071 12871 4075
rect 12807 4015 12811 4071
rect 12811 4015 12867 4071
rect 12867 4015 12871 4071
rect 12807 4011 12871 4015
rect 12887 4071 12951 4075
rect 12887 4015 12891 4071
rect 12891 4015 12947 4071
rect 12947 4015 12951 4071
rect 12887 4011 12951 4015
rect 12967 4071 13031 4075
rect 12967 4015 12971 4071
rect 12971 4015 13027 4071
rect 13027 4015 13031 4071
rect 12967 4011 13031 4015
rect 13047 4071 13111 4075
rect 13047 4015 13051 4071
rect 13051 4015 13107 4071
rect 13107 4015 13111 4071
rect 13047 4011 13111 4015
<< metal4 >>
rect -3536 22530 -2536 22592
rect -3536 21654 -3474 22530
rect -2598 21654 -2536 22530
rect -3536 -1526 -2536 21654
rect -2056 21050 -1056 21112
rect -2056 20174 -1994 21050
rect -1118 20174 -1056 21050
rect -2056 13384 -1056 20174
rect 5416 21066 6416 22592
rect 5416 20190 5478 21066
rect 6354 20190 6416 21066
rect -2056 12508 -1994 13384
rect -1118 12508 -1056 13384
rect -2056 -46 -1056 12508
rect -576 19570 424 19632
rect -576 18694 -514 19570
rect 362 18694 424 19570
rect -576 9593 424 18694
rect -576 8717 -514 9593
rect 362 8717 424 9593
rect -576 1434 424 8717
rect 904 18090 1904 18152
rect 904 17214 966 18090
rect 1842 17214 1904 18090
rect 904 2914 1904 17214
rect 904 2038 966 2914
rect 1842 2038 1904 2914
rect 904 1976 1904 2038
rect 5416 13400 6416 20190
rect 7440 22517 8197 22592
rect 7440 21641 7544 22517
rect 8100 21641 8197 22517
rect 7440 16237 8197 21641
rect 7440 16173 7451 16237
rect 7515 16173 7531 16237
rect 7595 16173 7611 16237
rect 7675 16173 7691 16237
rect 7755 16173 7817 16237
rect 7881 16173 7897 16237
rect 7961 16173 7977 16237
rect 8041 16173 8057 16237
rect 8121 16173 8197 16237
rect 7440 16118 8197 16173
rect 7440 16054 7451 16118
rect 7515 16054 7531 16118
rect 7595 16054 7611 16118
rect 7675 16054 7691 16118
rect 7755 16054 7817 16118
rect 7881 16054 7897 16118
rect 7961 16054 7977 16118
rect 8041 16054 8057 16118
rect 8121 16054 8197 16118
rect 7440 16042 8197 16054
rect 10170 18068 10927 22592
rect 10170 17192 10274 18068
rect 10830 17192 10927 18068
rect 10170 16237 10927 17192
rect 10170 16173 10181 16237
rect 10245 16173 10261 16237
rect 10325 16173 10341 16237
rect 10405 16173 10421 16237
rect 10485 16173 10547 16237
rect 10611 16173 10627 16237
rect 10691 16173 10707 16237
rect 10771 16173 10787 16237
rect 10851 16173 10927 16237
rect 10170 16118 10927 16173
rect 10170 16054 10181 16118
rect 10245 16054 10261 16118
rect 10325 16054 10341 16118
rect 10405 16054 10421 16118
rect 10485 16054 10547 16118
rect 10611 16054 10627 16118
rect 10691 16054 10707 16118
rect 10771 16054 10787 16118
rect 10851 16054 10927 16118
rect 10170 16042 10927 16054
rect 12130 19573 13130 22592
rect 20936 22530 21936 22592
rect 20936 21654 20998 22530
rect 21874 21654 21936 22530
rect 19456 21050 20456 21112
rect 19456 20174 19518 21050
rect 20394 20174 20456 21050
rect 12130 18697 12192 19573
rect 13068 18697 13130 19573
rect 5416 12524 5478 13400
rect 6354 12524 6416 13400
rect 5416 4187 6416 12524
rect 5416 4123 5427 4187
rect 5491 4123 5507 4187
rect 5571 4123 5587 4187
rect 5651 4123 5667 4187
rect 5731 4123 6093 4187
rect 6157 4123 6173 4187
rect 6237 4123 6253 4187
rect 6317 4123 6333 4187
rect 6397 4123 6416 4187
rect 5416 4068 6416 4123
rect 5416 4004 5427 4068
rect 5491 4004 5507 4068
rect 5571 4004 5587 4068
rect 5651 4004 5667 4068
rect 5731 4004 6093 4068
rect 6157 4004 6173 4068
rect 6237 4004 6253 4068
rect 6317 4004 6333 4068
rect 6397 4004 6416 4068
rect -576 558 -514 1434
rect 362 558 424 1434
rect -576 496 424 558
rect -2056 -922 -1994 -46
rect -1118 -922 -1056 -46
rect -2056 -984 -1056 -922
rect 5416 -56 6416 4004
rect 5416 -932 5478 -56
rect 6354 -932 6416 -56
rect -3536 -2402 -3474 -1526
rect -2598 -2402 -2536 -1526
rect -3536 -2464 -2536 -2402
rect 5416 -2464 6416 -932
rect 12130 9596 13130 18697
rect 17976 19570 18976 19632
rect 17976 18694 18038 19570
rect 18914 18694 18976 19570
rect 12130 8720 12192 9596
rect 13068 8720 13130 9596
rect 12130 4194 13130 8720
rect 12130 4130 12141 4194
rect 12205 4130 12221 4194
rect 12285 4130 12301 4194
rect 12365 4130 12381 4194
rect 12445 4130 12807 4194
rect 12871 4130 12887 4194
rect 12951 4130 12967 4194
rect 13031 4130 13047 4194
rect 13111 4130 13130 4194
rect 12130 4075 13130 4130
rect 12130 4011 12141 4075
rect 12205 4011 12221 4075
rect 12285 4011 12301 4075
rect 12365 4011 12381 4075
rect 12445 4011 12807 4075
rect 12871 4011 12887 4075
rect 12951 4011 12967 4075
rect 13031 4011 13047 4075
rect 13111 4011 13130 4075
rect 12130 1429 13130 4011
rect 16496 18090 17496 18152
rect 16496 17214 16558 18090
rect 17434 17214 17496 18090
rect 16496 2914 17496 17214
rect 16496 2038 16558 2914
rect 17434 2038 17496 2914
rect 16496 1976 17496 2038
rect 17976 9593 18976 18694
rect 17976 8717 18038 9593
rect 18914 8717 18976 9593
rect 12130 553 12192 1429
rect 13068 553 13130 1429
rect 12130 -2464 13130 553
rect 17976 1434 18976 8717
rect 17976 558 18038 1434
rect 18914 558 18976 1434
rect 17976 496 18976 558
rect 19456 13384 20456 20174
rect 19456 12508 19518 13384
rect 20394 12508 20456 13384
rect 19456 -46 20456 12508
rect 19456 -922 19518 -46
rect 20394 -922 20456 -46
rect 19456 -984 20456 -922
rect 20936 -1526 21936 21654
rect 20936 -2402 20998 -1526
rect 21874 -2402 21936 -1526
rect 20936 -2464 21936 -2402
<< via4 >>
rect -3474 21654 -2598 22530
rect -1994 20174 -1118 21050
rect 5478 20190 6354 21066
rect -1994 12508 -1118 13384
rect -514 18694 362 19570
rect -514 8717 362 9593
rect 966 17214 1842 18090
rect 966 2038 1842 2914
rect 7544 21641 8100 22517
rect 10274 17192 10830 18068
rect 20998 21654 21874 22530
rect 19518 20174 20394 21050
rect 12192 18697 13068 19573
rect 5478 12524 6354 13400
rect -514 558 362 1434
rect -1994 -922 -1118 -46
rect 5478 -932 6354 -56
rect -3474 -2402 -2598 -1526
rect 18038 18694 18914 19570
rect 12192 8720 13068 9596
rect 16558 17214 17434 18090
rect 16558 2038 17434 2914
rect 18038 8717 18914 9593
rect 12192 553 13068 1429
rect 18038 558 18914 1434
rect 19518 12508 20394 13384
rect 19518 -922 20394 -46
rect 20998 -2402 21874 -1526
<< metal5 >>
rect -3536 22530 21936 22592
rect -3536 21654 -3474 22530
rect -2598 22517 20998 22530
rect -2598 21654 7544 22517
rect -3536 21641 7544 21654
rect 8100 21654 20998 22517
rect 21874 21654 21936 22530
rect 8100 21641 21936 21654
rect -3536 21592 21936 21641
rect -2056 21066 20456 21112
rect -2056 21050 5478 21066
rect -2056 20174 -1994 21050
rect -1118 20190 5478 21050
rect 6354 21050 20456 21066
rect 6354 20190 19518 21050
rect -1118 20174 19518 20190
rect 20394 20174 20456 21050
rect -2056 20112 20456 20174
rect -576 19573 18976 19632
rect -576 19570 12192 19573
rect -576 18694 -514 19570
rect 362 18697 12192 19570
rect 13068 19570 18976 19573
rect 13068 18697 18038 19570
rect 362 18694 18038 18697
rect 18914 18694 18976 19570
rect -576 18632 18976 18694
rect 904 18090 17496 18152
rect 904 17214 966 18090
rect 1842 18068 16558 18090
rect 1842 17214 10274 18068
rect 904 17192 10274 17214
rect 10830 17214 16558 18068
rect 17434 17214 17496 18090
rect 10830 17192 17496 17214
rect 904 17152 17496 17192
rect -2056 13400 20456 13446
rect -2056 13384 5478 13400
rect -2056 12508 -1994 13384
rect -1118 12524 5478 13384
rect 6354 13384 20456 13400
rect 6354 12524 19518 13384
rect -1118 12508 19518 12524
rect 20394 12508 20456 13384
rect -2056 12446 20456 12508
rect -576 9596 18976 9655
rect -576 9593 12192 9596
rect -576 8717 -514 9593
rect 362 8720 12192 9593
rect 13068 9593 18976 9596
rect 13068 8720 18038 9593
rect 362 8717 18038 8720
rect 18914 8717 18976 9593
rect -576 8655 18976 8717
rect 904 2914 17496 2976
rect 904 2038 966 2914
rect 1842 2038 16558 2914
rect 17434 2038 17496 2914
rect 904 1976 17496 2038
rect -576 1434 18976 1496
rect -576 558 -514 1434
rect 362 1429 18038 1434
rect 362 558 12192 1429
rect -576 553 12192 558
rect 13068 558 18038 1429
rect 18914 558 18976 1434
rect 13068 553 18976 558
rect -576 496 18976 553
rect -2056 -46 20456 16
rect -2056 -922 -1994 -46
rect -1118 -56 19518 -46
rect -1118 -922 5478 -56
rect -2056 -932 5478 -922
rect 6354 -922 19518 -56
rect 20394 -922 20456 -46
rect 6354 -932 20456 -922
rect -2056 -984 20456 -932
rect -3536 -1526 21936 -1464
rect -3536 -2402 -3474 -1526
rect -2598 -2402 20998 -1526
rect 21874 -2402 21936 -1526
rect -3536 -2464 21936 -2402
use sky130_ef_ip__rc_osc_500k  mprj
timestamp 1527881472
transform 0 -1 14561 1 0 4000
box 0 0 12242 10724
<< labels >>
flabel metal2 s 9006 20076 9118 21516 0 FreeSans 560 90 0 0 dout
port 1 nsew
flabel metal2 s 9650 20076 9762 21516 0 FreeSans 560 90 0 0 ena
port 2 nsew
flabel metal4 s 5416 -2464 6416 22592 0 FreeSans 9600 90 0 0 vdda1
port 4 nsew
flabel metal4 s 12130 -2464 13130 22592 0 FreeSans 9600 90 0 0 vssa1
port 5 nsew
flabel metal4 s 16496 1976 17496 18152 0 FreeSans 9600 90 0 0 vccd1
port 3 nsew
flabel metal4 s 904 1976 1904 18152 0 FreeSans 9600 90 0 0 vccd1
port 3 nsew
flabel metal4 s 19456 -984 20456 21112 0 FreeSans 9600 90 0 0 vdda1
port 4 nsew
flabel metal4 s -2056 -984 -1056 21112 0 FreeSans 9600 90 0 0 vdda1
port 4 nsew
flabel metal4 s 17976 496 18976 19632 0 FreeSans 9600 90 0 0 vssa1
port 5 nsew
flabel metal4 s -576 496 424 19632 0 FreeSans 9600 90 0 0 vssa1
port 5 nsew
flabel metal4 s 20936 -2464 21936 22592 0 FreeSans 9600 90 0 0 vssd1
port 6 nsew
flabel metal4 s -3536 -2464 -2536 22592 0 FreeSans 9600 90 0 0 vssd1
port 6 nsew
flabel metal5 s -2056 12446 20456 13446 0 FreeSans 6400 0 0 0 vdda1
port 4 nsew
flabel metal5 s -576 8655 18976 9655 0 FreeSans 6400 0 0 0 vssa1
port 5 nsew
flabel metal5 s 904 17152 17496 18152 0 FreeSans 6400 0 0 0 vccd1
port 3 nsew
flabel metal5 s 904 1976 17496 2976 0 FreeSans 6400 0 0 0 vccd1
port 3 nsew
flabel metal5 s -2056 20112 20456 21112 0 FreeSans 6400 0 0 0 vdda1
port 4 nsew
flabel metal5 s -2056 -984 20456 16 0 FreeSans 6400 0 0 0 vdda1
port 4 nsew
flabel metal5 s -576 18632 18976 19632 0 FreeSans 6400 0 0 0 vssa1
port 5 nsew
flabel metal5 s -576 496 18976 1496 0 FreeSans 6400 0 0 0 vssa1
port 5 nsew
flabel metal5 s -3536 21592 21936 22592 0 FreeSans 6400 0 0 0 vssd1
port 6 nsew
flabel metal5 s -3536 -2464 21936 -1464 0 FreeSans 6400 0 0 0 vssd1
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 18412 20556
<< end >>

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__rc_osc_500k_DI
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__rc_osc_500k_DI ;
  ORIGIN 0.000 0.000 ;
  SIZE 54.360 BY 138.695 ;
  PIN dout
    ANTENNADIFFAREA 0.556800 ;
    PORT
      LAYER met2 ;
        RECT 26.445 137.015 27.005 144.215 ;
    END
  END dout
  PIN ena
    ANTENNAGATEAREA 0.858000 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 29.665 137.015 30.225 144.215 ;
    END
  END ena
  PIN vssd1
    ANTENNADIFFAREA 6.628900 ;
    PORT
      LAYER met4 ;
        RECT 18.615 92.530 21.715 138.695 ;
    END
  END vssd1
  PIN vccd1
    ANTENNADIFFAREA 4.280700 ;
    PORT
      LAYER met4 ;
        RECT 32.265 92.530 35.365 138.695 ;
    END
  END vccd1
  PIN vdda1
    ANTENNADIFFAREA 148.310989 ;
    PORT
      LAYER met4 ;
        RECT 8.495 0.000 13.495 138.695 ;
    END
  END vdda1
  PIN vssa1
    ANTENNADIFFAREA 114.014595 ;
    PORT
      LAYER met4 ;
        RECT 42.065 0.000 47.065 138.695 ;
    END
  END vssa1
  OBS
      LAYER nwell ;
        RECT 0.600 91.920 20.970 93.530 ;
        RECT 0.600 33.930 2.210 91.920 ;
        RECT 0.600 32.320 54.220 33.930 ;
      LAYER li1 ;
        RECT 1.040 32.750 53.755 93.075 ;
      LAYER met1 ;
        RECT 3.220 32.750 51.630 93.530 ;
      LAYER met2 ;
        RECT 5.740 136.735 26.165 138.215 ;
        RECT 27.285 136.735 29.385 138.215 ;
        RECT 30.505 136.735 48.880 138.215 ;
        RECT 5.740 32.320 48.880 136.735 ;
      LAYER met3 ;
        RECT 8.495 32.315 47.065 93.530 ;
      LAYER met4 ;
        RECT 26.230 43.875 36.370 69.655 ;
  END
END sky130_ef_ip__rc_osc_500k_DI
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1527949378
<< checkpaint >>
rect 2577 -3724 15821 24935
<< via1 >>
rect 7452 16183 7504 16235
rect 7516 16183 7568 16235
rect 7580 16183 7632 16235
rect 7644 16183 7696 16235
rect 7820 16183 7872 16235
rect 7884 16183 7936 16235
rect 7948 16183 8000 16235
rect 8126 16182 8178 16234
rect 10186 16183 10238 16235
rect 10250 16183 10302 16235
rect 10314 16183 10366 16235
rect 10378 16183 10430 16235
rect 10554 16183 10606 16235
rect 10618 16183 10670 16235
rect 10682 16183 10734 16235
rect 10860 16182 10912 16234
rect 7452 16093 7504 16145
rect 7516 16093 7568 16145
rect 7580 16093 7632 16145
rect 7644 16093 7696 16145
rect 7820 16093 7872 16145
rect 7884 16093 7936 16145
rect 7948 16093 8000 16145
rect 8126 16092 8178 16144
rect 10186 16093 10238 16145
rect 10250 16093 10302 16145
rect 10314 16093 10366 16145
rect 10378 16093 10430 16145
rect 10554 16093 10606 16145
rect 10618 16093 10670 16145
rect 10682 16093 10734 16145
rect 10860 16092 10912 16144
<< metal2 >>
rect 9006 20210 9118 21516
rect 9650 20316 9762 21516
rect 8864 20182 9118 20210
rect 7440 16235 8197 16242
rect 7440 16183 7452 16235
rect 7504 16233 7516 16235
rect 7568 16233 7580 16235
rect 7632 16233 7644 16235
rect 7696 16233 7820 16235
rect 7872 16233 7884 16235
rect 7936 16233 7948 16235
rect 8000 16234 8197 16235
rect 8000 16233 8126 16234
rect 7511 16183 7516 16233
rect 7751 16183 7820 16233
rect 7877 16183 7884 16233
rect 7440 16177 7455 16183
rect 7511 16177 7535 16183
rect 7591 16177 7615 16183
rect 7671 16177 7695 16183
rect 7751 16177 7821 16183
rect 7877 16177 7901 16183
rect 7957 16177 7981 16183
rect 8037 16177 8061 16233
rect 8117 16182 8126 16233
rect 8178 16182 8197 16234
rect 8117 16177 8197 16182
rect 7440 16145 8197 16177
rect 7440 16093 7452 16145
rect 7504 16114 7516 16145
rect 7568 16114 7580 16145
rect 7632 16114 7644 16145
rect 7696 16114 7820 16145
rect 7872 16114 7884 16145
rect 7936 16114 7948 16145
rect 8000 16144 8197 16145
rect 8000 16114 8126 16144
rect 7511 16093 7516 16114
rect 7751 16093 7820 16114
rect 7877 16093 7884 16114
rect 7440 16058 7455 16093
rect 7511 16058 7535 16093
rect 7591 16058 7615 16093
rect 7671 16058 7695 16093
rect 7751 16058 7821 16093
rect 7877 16058 7901 16093
rect 7957 16058 7981 16093
rect 8037 16058 8061 16114
rect 8117 16092 8126 16114
rect 8178 16092 8197 16144
rect 8864 16116 8892 20182
rect 9006 20076 9118 20182
rect 9641 20076 9762 20316
rect 9641 20074 9669 20076
rect 9600 20046 9669 20074
rect 9600 16116 9628 20046
rect 10170 16235 10927 16242
rect 10170 16233 10186 16235
rect 10238 16233 10250 16235
rect 10302 16233 10314 16235
rect 10366 16233 10378 16235
rect 10430 16233 10554 16235
rect 10606 16233 10618 16235
rect 10670 16233 10682 16235
rect 10734 16234 10927 16235
rect 10734 16233 10860 16234
rect 10170 16177 10185 16233
rect 10241 16183 10250 16233
rect 10241 16177 10265 16183
rect 10321 16177 10345 16183
rect 10401 16177 10425 16183
rect 10481 16177 10551 16233
rect 10607 16183 10618 16233
rect 10607 16177 10631 16183
rect 10687 16177 10711 16183
rect 10767 16177 10791 16233
rect 10847 16182 10860 16233
rect 10912 16182 10927 16234
rect 10847 16177 10927 16182
rect 10170 16145 10927 16177
rect 8117 16058 8197 16092
rect 7440 16042 8197 16058
rect 10170 16114 10186 16145
rect 10238 16114 10250 16145
rect 10302 16114 10314 16145
rect 10366 16114 10378 16145
rect 10430 16114 10554 16145
rect 10606 16114 10618 16145
rect 10670 16114 10682 16145
rect 10734 16144 10927 16145
rect 10734 16114 10860 16144
rect 10170 16058 10185 16114
rect 10241 16093 10250 16114
rect 10241 16058 10265 16093
rect 10321 16058 10345 16093
rect 10401 16058 10425 16093
rect 10481 16058 10551 16114
rect 10607 16093 10618 16114
rect 10607 16058 10631 16093
rect 10687 16058 10711 16093
rect 10767 16058 10791 16114
rect 10847 16092 10860 16114
rect 10912 16092 10927 16144
rect 10847 16058 10927 16092
rect 10170 16042 10927 16058
<< via2 >>
rect 7455 16183 7504 16233
rect 7504 16183 7511 16233
rect 7535 16183 7568 16233
rect 7568 16183 7580 16233
rect 7580 16183 7591 16233
rect 7615 16183 7632 16233
rect 7632 16183 7644 16233
rect 7644 16183 7671 16233
rect 7695 16183 7696 16233
rect 7696 16183 7751 16233
rect 7821 16183 7872 16233
rect 7872 16183 7877 16233
rect 7901 16183 7936 16233
rect 7936 16183 7948 16233
rect 7948 16183 7957 16233
rect 7981 16183 8000 16233
rect 8000 16183 8037 16233
rect 7455 16177 7511 16183
rect 7535 16177 7591 16183
rect 7615 16177 7671 16183
rect 7695 16177 7751 16183
rect 7821 16177 7877 16183
rect 7901 16177 7957 16183
rect 7981 16177 8037 16183
rect 8061 16177 8117 16233
rect 7455 16093 7504 16114
rect 7504 16093 7511 16114
rect 7535 16093 7568 16114
rect 7568 16093 7580 16114
rect 7580 16093 7591 16114
rect 7615 16093 7632 16114
rect 7632 16093 7644 16114
rect 7644 16093 7671 16114
rect 7695 16093 7696 16114
rect 7696 16093 7751 16114
rect 7821 16093 7872 16114
rect 7872 16093 7877 16114
rect 7901 16093 7936 16114
rect 7936 16093 7948 16114
rect 7948 16093 7957 16114
rect 7981 16093 8000 16114
rect 8000 16093 8037 16114
rect 7455 16058 7511 16093
rect 7535 16058 7591 16093
rect 7615 16058 7671 16093
rect 7695 16058 7751 16093
rect 7821 16058 7877 16093
rect 7901 16058 7957 16093
rect 7981 16058 8037 16093
rect 8061 16058 8117 16114
rect 10185 16183 10186 16233
rect 10186 16183 10238 16233
rect 10238 16183 10241 16233
rect 10265 16183 10302 16233
rect 10302 16183 10314 16233
rect 10314 16183 10321 16233
rect 10345 16183 10366 16233
rect 10366 16183 10378 16233
rect 10378 16183 10401 16233
rect 10425 16183 10430 16233
rect 10430 16183 10481 16233
rect 10185 16177 10241 16183
rect 10265 16177 10321 16183
rect 10345 16177 10401 16183
rect 10425 16177 10481 16183
rect 10551 16183 10554 16233
rect 10554 16183 10606 16233
rect 10606 16183 10607 16233
rect 10631 16183 10670 16233
rect 10670 16183 10682 16233
rect 10682 16183 10687 16233
rect 10711 16183 10734 16233
rect 10734 16183 10767 16233
rect 10551 16177 10607 16183
rect 10631 16177 10687 16183
rect 10711 16177 10767 16183
rect 10791 16177 10847 16233
rect 10185 16093 10186 16114
rect 10186 16093 10238 16114
rect 10238 16093 10241 16114
rect 10265 16093 10302 16114
rect 10302 16093 10314 16114
rect 10314 16093 10321 16114
rect 10345 16093 10366 16114
rect 10366 16093 10378 16114
rect 10378 16093 10401 16114
rect 10425 16093 10430 16114
rect 10430 16093 10481 16114
rect 10185 16058 10241 16093
rect 10265 16058 10321 16093
rect 10345 16058 10401 16093
rect 10425 16058 10481 16093
rect 10551 16093 10554 16114
rect 10554 16093 10606 16114
rect 10606 16093 10607 16114
rect 10631 16093 10670 16114
rect 10670 16093 10682 16114
rect 10682 16093 10687 16114
rect 10711 16093 10734 16114
rect 10734 16093 10767 16114
rect 10551 16058 10607 16093
rect 10631 16058 10687 16093
rect 10711 16058 10767 16093
rect 10791 16058 10847 16114
rect 5431 15947 5487 16003
rect 5511 15947 5567 16003
rect 5591 15947 5647 16003
rect 5671 15947 5727 16003
rect 6097 15947 6153 16003
rect 6177 15947 6233 16003
rect 6257 15947 6313 16003
rect 6337 15947 6393 16003
rect 12145 15974 12201 16030
rect 12225 15974 12281 16030
rect 12305 15974 12361 16030
rect 12385 15974 12441 16030
rect 12811 15974 12867 16030
rect 12891 15974 12947 16030
rect 12971 15974 13027 16030
rect 13051 15974 13107 16030
rect 5431 15828 5487 15884
rect 5511 15828 5567 15884
rect 5591 15828 5647 15884
rect 5671 15828 5727 15884
rect 6097 15828 6153 15884
rect 6177 15828 6233 15884
rect 6257 15828 6313 15884
rect 6337 15828 6393 15884
rect 12145 15855 12201 15911
rect 12225 15855 12281 15911
rect 12305 15855 12361 15911
rect 12385 15855 12441 15911
rect 12811 15855 12867 15911
rect 12891 15855 12947 15911
rect 12971 15855 13027 15911
rect 13051 15855 13107 15911
rect 5431 4127 5487 4183
rect 5511 4127 5567 4183
rect 5591 4127 5647 4183
rect 5671 4127 5727 4183
rect 6097 4127 6153 4183
rect 6177 4127 6233 4183
rect 6257 4127 6313 4183
rect 6337 4127 6393 4183
rect 12145 4134 12201 4190
rect 12225 4134 12281 4190
rect 12305 4134 12361 4190
rect 12385 4134 12441 4190
rect 12811 4134 12867 4190
rect 12891 4134 12947 4190
rect 12971 4134 13027 4190
rect 13051 4134 13107 4190
rect 5431 4008 5487 4064
rect 5511 4008 5567 4064
rect 5591 4008 5647 4064
rect 5671 4008 5727 4064
rect 6097 4008 6153 4064
rect 6177 4008 6233 4064
rect 6257 4008 6313 4064
rect 6337 4008 6393 4064
rect 12145 4015 12201 4071
rect 12225 4015 12281 4071
rect 12305 4015 12361 4071
rect 12385 4015 12441 4071
rect 12811 4015 12867 4071
rect 12891 4015 12947 4071
rect 12971 4015 13027 4071
rect 13051 4015 13107 4071
<< metal3 >>
rect 7440 16237 8197 16242
rect 7440 16173 7451 16237
rect 7515 16173 7531 16237
rect 7595 16173 7611 16237
rect 7675 16173 7691 16237
rect 7755 16173 7817 16237
rect 7881 16173 7897 16237
rect 7961 16173 7977 16237
rect 8041 16173 8057 16237
rect 8121 16173 8197 16237
rect 5416 16007 6416 16161
rect 7440 16118 8197 16173
rect 7440 16054 7451 16118
rect 7515 16054 7531 16118
rect 7595 16054 7611 16118
rect 7675 16054 7691 16118
rect 7755 16054 7817 16118
rect 7881 16054 7897 16118
rect 7961 16054 7977 16118
rect 8041 16054 8057 16118
rect 8121 16054 8197 16118
rect 7440 16042 8197 16054
rect 10170 16237 10927 16242
rect 10170 16173 10181 16237
rect 10245 16173 10261 16237
rect 10325 16173 10341 16237
rect 10405 16173 10421 16237
rect 10485 16173 10547 16237
rect 10611 16173 10627 16237
rect 10691 16173 10707 16237
rect 10771 16173 10787 16237
rect 10851 16173 10927 16237
rect 10170 16118 10927 16173
rect 10170 16054 10181 16118
rect 10245 16054 10261 16118
rect 10325 16054 10341 16118
rect 10405 16054 10421 16118
rect 10485 16054 10547 16118
rect 10611 16054 10627 16118
rect 10691 16054 10707 16118
rect 10771 16054 10787 16118
rect 10851 16054 10927 16118
rect 10170 16042 10927 16054
rect 5416 15943 5427 16007
rect 5491 15943 5507 16007
rect 5571 15943 5587 16007
rect 5651 15943 5667 16007
rect 5731 15943 6093 16007
rect 6157 15943 6173 16007
rect 6237 15943 6253 16007
rect 6317 15943 6333 16007
rect 6397 15943 6416 16007
rect 5416 15888 6416 15943
rect 5416 15824 5427 15888
rect 5491 15824 5507 15888
rect 5571 15824 5587 15888
rect 5651 15824 5667 15888
rect 5731 15824 6093 15888
rect 6157 15824 6173 15888
rect 6237 15824 6253 15888
rect 6317 15824 6333 15888
rect 6397 15824 6416 15888
rect 12130 16034 13130 16181
rect 12130 15970 12141 16034
rect 12205 15970 12221 16034
rect 12285 15970 12301 16034
rect 12365 15970 12381 16034
rect 12445 15970 12807 16034
rect 12871 15970 12887 16034
rect 12951 15970 12967 16034
rect 13031 15970 13047 16034
rect 13111 15970 13130 16034
rect 12130 15915 13130 15970
rect 12130 15851 12141 15915
rect 12205 15851 12221 15915
rect 12285 15851 12301 15915
rect 12365 15851 12381 15915
rect 12445 15851 12807 15915
rect 12871 15851 12887 15915
rect 12951 15851 12967 15915
rect 13031 15851 13047 15915
rect 13111 15851 13130 15915
rect 12130 15839 13130 15851
rect 5416 15819 6416 15824
rect 5416 4187 6416 4341
rect 5416 4123 5427 4187
rect 5491 4123 5507 4187
rect 5571 4123 5587 4187
rect 5651 4123 5667 4187
rect 5731 4123 6093 4187
rect 6157 4123 6173 4187
rect 6237 4123 6253 4187
rect 6317 4123 6333 4187
rect 6397 4123 6416 4187
rect 5416 4068 6416 4123
rect 5416 4004 5427 4068
rect 5491 4004 5507 4068
rect 5571 4004 5587 4068
rect 5651 4004 5667 4068
rect 5731 4004 6093 4068
rect 6157 4004 6173 4068
rect 6237 4004 6253 4068
rect 6317 4004 6333 4068
rect 6397 4004 6416 4068
rect 5416 3999 6416 4004
rect 12130 4194 13130 4341
rect 12130 4130 12141 4194
rect 12205 4130 12221 4194
rect 12285 4130 12301 4194
rect 12365 4130 12381 4194
rect 12445 4130 12807 4194
rect 12871 4130 12887 4194
rect 12951 4130 12967 4194
rect 13031 4130 13047 4194
rect 13111 4130 13130 4194
rect 12130 4075 13130 4130
rect 12130 4011 12141 4075
rect 12205 4011 12221 4075
rect 12285 4011 12301 4075
rect 12365 4011 12381 4075
rect 12445 4011 12807 4075
rect 12871 4011 12887 4075
rect 12951 4011 12967 4075
rect 13031 4011 13047 4075
rect 13111 4011 13130 4075
rect 12130 3999 13130 4011
<< via3 >>
rect 7451 16233 7515 16237
rect 7451 16177 7455 16233
rect 7455 16177 7511 16233
rect 7511 16177 7515 16233
rect 7451 16173 7515 16177
rect 7531 16233 7595 16237
rect 7531 16177 7535 16233
rect 7535 16177 7591 16233
rect 7591 16177 7595 16233
rect 7531 16173 7595 16177
rect 7611 16233 7675 16237
rect 7611 16177 7615 16233
rect 7615 16177 7671 16233
rect 7671 16177 7675 16233
rect 7611 16173 7675 16177
rect 7691 16233 7755 16237
rect 7691 16177 7695 16233
rect 7695 16177 7751 16233
rect 7751 16177 7755 16233
rect 7691 16173 7755 16177
rect 7817 16233 7881 16237
rect 7817 16177 7821 16233
rect 7821 16177 7877 16233
rect 7877 16177 7881 16233
rect 7817 16173 7881 16177
rect 7897 16233 7961 16237
rect 7897 16177 7901 16233
rect 7901 16177 7957 16233
rect 7957 16177 7961 16233
rect 7897 16173 7961 16177
rect 7977 16233 8041 16237
rect 7977 16177 7981 16233
rect 7981 16177 8037 16233
rect 8037 16177 8041 16233
rect 7977 16173 8041 16177
rect 8057 16233 8121 16237
rect 8057 16177 8061 16233
rect 8061 16177 8117 16233
rect 8117 16177 8121 16233
rect 8057 16173 8121 16177
rect 7451 16114 7515 16118
rect 7451 16058 7455 16114
rect 7455 16058 7511 16114
rect 7511 16058 7515 16114
rect 7451 16054 7515 16058
rect 7531 16114 7595 16118
rect 7531 16058 7535 16114
rect 7535 16058 7591 16114
rect 7591 16058 7595 16114
rect 7531 16054 7595 16058
rect 7611 16114 7675 16118
rect 7611 16058 7615 16114
rect 7615 16058 7671 16114
rect 7671 16058 7675 16114
rect 7611 16054 7675 16058
rect 7691 16114 7755 16118
rect 7691 16058 7695 16114
rect 7695 16058 7751 16114
rect 7751 16058 7755 16114
rect 7691 16054 7755 16058
rect 7817 16114 7881 16118
rect 7817 16058 7821 16114
rect 7821 16058 7877 16114
rect 7877 16058 7881 16114
rect 7817 16054 7881 16058
rect 7897 16114 7961 16118
rect 7897 16058 7901 16114
rect 7901 16058 7957 16114
rect 7957 16058 7961 16114
rect 7897 16054 7961 16058
rect 7977 16114 8041 16118
rect 7977 16058 7981 16114
rect 7981 16058 8037 16114
rect 8037 16058 8041 16114
rect 7977 16054 8041 16058
rect 8057 16114 8121 16118
rect 8057 16058 8061 16114
rect 8061 16058 8117 16114
rect 8117 16058 8121 16114
rect 8057 16054 8121 16058
rect 10181 16233 10245 16237
rect 10181 16177 10185 16233
rect 10185 16177 10241 16233
rect 10241 16177 10245 16233
rect 10181 16173 10245 16177
rect 10261 16233 10325 16237
rect 10261 16177 10265 16233
rect 10265 16177 10321 16233
rect 10321 16177 10325 16233
rect 10261 16173 10325 16177
rect 10341 16233 10405 16237
rect 10341 16177 10345 16233
rect 10345 16177 10401 16233
rect 10401 16177 10405 16233
rect 10341 16173 10405 16177
rect 10421 16233 10485 16237
rect 10421 16177 10425 16233
rect 10425 16177 10481 16233
rect 10481 16177 10485 16233
rect 10421 16173 10485 16177
rect 10547 16233 10611 16237
rect 10547 16177 10551 16233
rect 10551 16177 10607 16233
rect 10607 16177 10611 16233
rect 10547 16173 10611 16177
rect 10627 16233 10691 16237
rect 10627 16177 10631 16233
rect 10631 16177 10687 16233
rect 10687 16177 10691 16233
rect 10627 16173 10691 16177
rect 10707 16233 10771 16237
rect 10707 16177 10711 16233
rect 10711 16177 10767 16233
rect 10767 16177 10771 16233
rect 10707 16173 10771 16177
rect 10787 16233 10851 16237
rect 10787 16177 10791 16233
rect 10791 16177 10847 16233
rect 10847 16177 10851 16233
rect 10787 16173 10851 16177
rect 10181 16114 10245 16118
rect 10181 16058 10185 16114
rect 10185 16058 10241 16114
rect 10241 16058 10245 16114
rect 10181 16054 10245 16058
rect 10261 16114 10325 16118
rect 10261 16058 10265 16114
rect 10265 16058 10321 16114
rect 10321 16058 10325 16114
rect 10261 16054 10325 16058
rect 10341 16114 10405 16118
rect 10341 16058 10345 16114
rect 10345 16058 10401 16114
rect 10401 16058 10405 16114
rect 10341 16054 10405 16058
rect 10421 16114 10485 16118
rect 10421 16058 10425 16114
rect 10425 16058 10481 16114
rect 10481 16058 10485 16114
rect 10421 16054 10485 16058
rect 10547 16114 10611 16118
rect 10547 16058 10551 16114
rect 10551 16058 10607 16114
rect 10607 16058 10611 16114
rect 10547 16054 10611 16058
rect 10627 16114 10691 16118
rect 10627 16058 10631 16114
rect 10631 16058 10687 16114
rect 10687 16058 10691 16114
rect 10627 16054 10691 16058
rect 10707 16114 10771 16118
rect 10707 16058 10711 16114
rect 10711 16058 10767 16114
rect 10767 16058 10771 16114
rect 10707 16054 10771 16058
rect 10787 16114 10851 16118
rect 10787 16058 10791 16114
rect 10791 16058 10847 16114
rect 10847 16058 10851 16114
rect 10787 16054 10851 16058
rect 5427 16003 5491 16007
rect 5427 15947 5431 16003
rect 5431 15947 5487 16003
rect 5487 15947 5491 16003
rect 5427 15943 5491 15947
rect 5507 16003 5571 16007
rect 5507 15947 5511 16003
rect 5511 15947 5567 16003
rect 5567 15947 5571 16003
rect 5507 15943 5571 15947
rect 5587 16003 5651 16007
rect 5587 15947 5591 16003
rect 5591 15947 5647 16003
rect 5647 15947 5651 16003
rect 5587 15943 5651 15947
rect 5667 16003 5731 16007
rect 5667 15947 5671 16003
rect 5671 15947 5727 16003
rect 5727 15947 5731 16003
rect 5667 15943 5731 15947
rect 6093 16003 6157 16007
rect 6093 15947 6097 16003
rect 6097 15947 6153 16003
rect 6153 15947 6157 16003
rect 6093 15943 6157 15947
rect 6173 16003 6237 16007
rect 6173 15947 6177 16003
rect 6177 15947 6233 16003
rect 6233 15947 6237 16003
rect 6173 15943 6237 15947
rect 6253 16003 6317 16007
rect 6253 15947 6257 16003
rect 6257 15947 6313 16003
rect 6313 15947 6317 16003
rect 6253 15943 6317 15947
rect 6333 16003 6397 16007
rect 6333 15947 6337 16003
rect 6337 15947 6393 16003
rect 6393 15947 6397 16003
rect 6333 15943 6397 15947
rect 5427 15884 5491 15888
rect 5427 15828 5431 15884
rect 5431 15828 5487 15884
rect 5487 15828 5491 15884
rect 5427 15824 5491 15828
rect 5507 15884 5571 15888
rect 5507 15828 5511 15884
rect 5511 15828 5567 15884
rect 5567 15828 5571 15884
rect 5507 15824 5571 15828
rect 5587 15884 5651 15888
rect 5587 15828 5591 15884
rect 5591 15828 5647 15884
rect 5647 15828 5651 15884
rect 5587 15824 5651 15828
rect 5667 15884 5731 15888
rect 5667 15828 5671 15884
rect 5671 15828 5727 15884
rect 5727 15828 5731 15884
rect 5667 15824 5731 15828
rect 6093 15884 6157 15888
rect 6093 15828 6097 15884
rect 6097 15828 6153 15884
rect 6153 15828 6157 15884
rect 6093 15824 6157 15828
rect 6173 15884 6237 15888
rect 6173 15828 6177 15884
rect 6177 15828 6233 15884
rect 6233 15828 6237 15884
rect 6173 15824 6237 15828
rect 6253 15884 6317 15888
rect 6253 15828 6257 15884
rect 6257 15828 6313 15884
rect 6313 15828 6317 15884
rect 6253 15824 6317 15828
rect 6333 15884 6397 15888
rect 6333 15828 6337 15884
rect 6337 15828 6393 15884
rect 6393 15828 6397 15884
rect 6333 15824 6397 15828
rect 12141 16030 12205 16034
rect 12141 15974 12145 16030
rect 12145 15974 12201 16030
rect 12201 15974 12205 16030
rect 12141 15970 12205 15974
rect 12221 16030 12285 16034
rect 12221 15974 12225 16030
rect 12225 15974 12281 16030
rect 12281 15974 12285 16030
rect 12221 15970 12285 15974
rect 12301 16030 12365 16034
rect 12301 15974 12305 16030
rect 12305 15974 12361 16030
rect 12361 15974 12365 16030
rect 12301 15970 12365 15974
rect 12381 16030 12445 16034
rect 12381 15974 12385 16030
rect 12385 15974 12441 16030
rect 12441 15974 12445 16030
rect 12381 15970 12445 15974
rect 12807 16030 12871 16034
rect 12807 15974 12811 16030
rect 12811 15974 12867 16030
rect 12867 15974 12871 16030
rect 12807 15970 12871 15974
rect 12887 16030 12951 16034
rect 12887 15974 12891 16030
rect 12891 15974 12947 16030
rect 12947 15974 12951 16030
rect 12887 15970 12951 15974
rect 12967 16030 13031 16034
rect 12967 15974 12971 16030
rect 12971 15974 13027 16030
rect 13027 15974 13031 16030
rect 12967 15970 13031 15974
rect 13047 16030 13111 16034
rect 13047 15974 13051 16030
rect 13051 15974 13107 16030
rect 13107 15974 13111 16030
rect 13047 15970 13111 15974
rect 12141 15911 12205 15915
rect 12141 15855 12145 15911
rect 12145 15855 12201 15911
rect 12201 15855 12205 15911
rect 12141 15851 12205 15855
rect 12221 15911 12285 15915
rect 12221 15855 12225 15911
rect 12225 15855 12281 15911
rect 12281 15855 12285 15911
rect 12221 15851 12285 15855
rect 12301 15911 12365 15915
rect 12301 15855 12305 15911
rect 12305 15855 12361 15911
rect 12361 15855 12365 15911
rect 12301 15851 12365 15855
rect 12381 15911 12445 15915
rect 12381 15855 12385 15911
rect 12385 15855 12441 15911
rect 12441 15855 12445 15911
rect 12381 15851 12445 15855
rect 12807 15911 12871 15915
rect 12807 15855 12811 15911
rect 12811 15855 12867 15911
rect 12867 15855 12871 15911
rect 12807 15851 12871 15855
rect 12887 15911 12951 15915
rect 12887 15855 12891 15911
rect 12891 15855 12947 15911
rect 12947 15855 12951 15911
rect 12887 15851 12951 15855
rect 12967 15911 13031 15915
rect 12967 15855 12971 15911
rect 12971 15855 13027 15911
rect 13027 15855 13031 15911
rect 12967 15851 13031 15855
rect 13047 15911 13111 15915
rect 13047 15855 13051 15911
rect 13051 15855 13107 15911
rect 13107 15855 13111 15911
rect 13047 15851 13111 15855
rect 5427 4183 5491 4187
rect 5427 4127 5431 4183
rect 5431 4127 5487 4183
rect 5487 4127 5491 4183
rect 5427 4123 5491 4127
rect 5507 4183 5571 4187
rect 5507 4127 5511 4183
rect 5511 4127 5567 4183
rect 5567 4127 5571 4183
rect 5507 4123 5571 4127
rect 5587 4183 5651 4187
rect 5587 4127 5591 4183
rect 5591 4127 5647 4183
rect 5647 4127 5651 4183
rect 5587 4123 5651 4127
rect 5667 4183 5731 4187
rect 5667 4127 5671 4183
rect 5671 4127 5727 4183
rect 5727 4127 5731 4183
rect 5667 4123 5731 4127
rect 6093 4183 6157 4187
rect 6093 4127 6097 4183
rect 6097 4127 6153 4183
rect 6153 4127 6157 4183
rect 6093 4123 6157 4127
rect 6173 4183 6237 4187
rect 6173 4127 6177 4183
rect 6177 4127 6233 4183
rect 6233 4127 6237 4183
rect 6173 4123 6237 4127
rect 6253 4183 6317 4187
rect 6253 4127 6257 4183
rect 6257 4127 6313 4183
rect 6313 4127 6317 4183
rect 6253 4123 6317 4127
rect 6333 4183 6397 4187
rect 6333 4127 6337 4183
rect 6337 4127 6393 4183
rect 6393 4127 6397 4183
rect 6333 4123 6397 4127
rect 5427 4064 5491 4068
rect 5427 4008 5431 4064
rect 5431 4008 5487 4064
rect 5487 4008 5491 4064
rect 5427 4004 5491 4008
rect 5507 4064 5571 4068
rect 5507 4008 5511 4064
rect 5511 4008 5567 4064
rect 5567 4008 5571 4064
rect 5507 4004 5571 4008
rect 5587 4064 5651 4068
rect 5587 4008 5591 4064
rect 5591 4008 5647 4064
rect 5647 4008 5651 4064
rect 5587 4004 5651 4008
rect 5667 4064 5731 4068
rect 5667 4008 5671 4064
rect 5671 4008 5727 4064
rect 5727 4008 5731 4064
rect 5667 4004 5731 4008
rect 6093 4064 6157 4068
rect 6093 4008 6097 4064
rect 6097 4008 6153 4064
rect 6153 4008 6157 4064
rect 6093 4004 6157 4008
rect 6173 4064 6237 4068
rect 6173 4008 6177 4064
rect 6177 4008 6233 4064
rect 6233 4008 6237 4064
rect 6173 4004 6237 4008
rect 6253 4064 6317 4068
rect 6253 4008 6257 4064
rect 6257 4008 6313 4064
rect 6313 4008 6317 4064
rect 6253 4004 6317 4008
rect 6333 4064 6397 4068
rect 6333 4008 6337 4064
rect 6337 4008 6393 4064
rect 6393 4008 6397 4064
rect 6333 4004 6397 4008
rect 12141 4190 12205 4194
rect 12141 4134 12145 4190
rect 12145 4134 12201 4190
rect 12201 4134 12205 4190
rect 12141 4130 12205 4134
rect 12221 4190 12285 4194
rect 12221 4134 12225 4190
rect 12225 4134 12281 4190
rect 12281 4134 12285 4190
rect 12221 4130 12285 4134
rect 12301 4190 12365 4194
rect 12301 4134 12305 4190
rect 12305 4134 12361 4190
rect 12361 4134 12365 4190
rect 12301 4130 12365 4134
rect 12381 4190 12445 4194
rect 12381 4134 12385 4190
rect 12385 4134 12441 4190
rect 12441 4134 12445 4190
rect 12381 4130 12445 4134
rect 12807 4190 12871 4194
rect 12807 4134 12811 4190
rect 12811 4134 12867 4190
rect 12867 4134 12871 4190
rect 12807 4130 12871 4134
rect 12887 4190 12951 4194
rect 12887 4134 12891 4190
rect 12891 4134 12947 4190
rect 12947 4134 12951 4190
rect 12887 4130 12951 4134
rect 12967 4190 13031 4194
rect 12967 4134 12971 4190
rect 12971 4134 13027 4190
rect 13027 4134 13031 4190
rect 12967 4130 13031 4134
rect 13047 4190 13111 4194
rect 13047 4134 13051 4190
rect 13051 4134 13107 4190
rect 13107 4134 13111 4190
rect 13047 4130 13111 4134
rect 12141 4071 12205 4075
rect 12141 4015 12145 4071
rect 12145 4015 12201 4071
rect 12201 4015 12205 4071
rect 12141 4011 12205 4015
rect 12221 4071 12285 4075
rect 12221 4015 12225 4071
rect 12225 4015 12281 4071
rect 12281 4015 12285 4071
rect 12221 4011 12285 4015
rect 12301 4071 12365 4075
rect 12301 4015 12305 4071
rect 12305 4015 12361 4071
rect 12361 4015 12365 4071
rect 12301 4011 12365 4015
rect 12381 4071 12445 4075
rect 12381 4015 12385 4071
rect 12385 4015 12441 4071
rect 12441 4015 12445 4071
rect 12381 4011 12445 4015
rect 12807 4071 12871 4075
rect 12807 4015 12811 4071
rect 12811 4015 12867 4071
rect 12867 4015 12871 4071
rect 12807 4011 12871 4015
rect 12887 4071 12951 4075
rect 12887 4015 12891 4071
rect 12891 4015 12947 4071
rect 12947 4015 12951 4071
rect 12887 4011 12951 4015
rect 12967 4071 13031 4075
rect 12967 4015 12971 4071
rect 12971 4015 13027 4071
rect 13027 4015 13031 4071
rect 12967 4011 13031 4015
rect 13047 4071 13111 4075
rect 13047 4015 13051 4071
rect 13051 4015 13107 4071
rect 13107 4015 13111 4071
rect 13047 4011 13111 4015
<< metal4 >>
rect 5416 16007 6416 22592
rect 7440 16237 8197 23675
rect 7440 16173 7451 16237
rect 7515 16173 7531 16237
rect 7595 16173 7611 16237
rect 7675 16173 7691 16237
rect 7755 16173 7817 16237
rect 7881 16173 7897 16237
rect 7961 16173 7977 16237
rect 8041 16173 8057 16237
rect 8121 16173 8197 16237
rect 7440 16118 8197 16173
rect 7440 16054 7451 16118
rect 7515 16054 7531 16118
rect 7595 16054 7611 16118
rect 7675 16054 7691 16118
rect 7755 16054 7817 16118
rect 7881 16054 7897 16118
rect 7961 16054 7977 16118
rect 8041 16054 8057 16118
rect 8121 16054 8197 16118
rect 7440 16042 8197 16054
rect 10170 16237 10927 23675
rect 10170 16173 10181 16237
rect 10245 16173 10261 16237
rect 10325 16173 10341 16237
rect 10405 16173 10421 16237
rect 10485 16173 10547 16237
rect 10611 16173 10627 16237
rect 10691 16173 10707 16237
rect 10771 16173 10787 16237
rect 10851 16173 10927 16237
rect 10170 16118 10927 16173
rect 10170 16054 10181 16118
rect 10245 16054 10261 16118
rect 10325 16054 10341 16118
rect 10405 16054 10421 16118
rect 10485 16054 10547 16118
rect 10611 16054 10627 16118
rect 10691 16054 10707 16118
rect 10771 16054 10787 16118
rect 10851 16054 10927 16118
rect 10170 16042 10927 16054
rect 5416 15943 5427 16007
rect 5491 15943 5507 16007
rect 5571 15943 5587 16007
rect 5651 15943 5667 16007
rect 5731 15943 6093 16007
rect 6157 15943 6173 16007
rect 6237 15943 6253 16007
rect 6317 15943 6333 16007
rect 6397 15943 6416 16007
rect 5416 15888 6416 15943
rect 5416 15824 5427 15888
rect 5491 15824 5507 15888
rect 5571 15824 5587 15888
rect 5651 15824 5667 15888
rect 5731 15824 6093 15888
rect 6157 15824 6173 15888
rect 6237 15824 6253 15888
rect 6317 15824 6333 15888
rect 6397 15824 6416 15888
rect 5416 4187 6416 15824
rect 5416 4123 5427 4187
rect 5491 4123 5507 4187
rect 5571 4123 5587 4187
rect 5651 4123 5667 4187
rect 5731 4123 6093 4187
rect 6157 4123 6173 4187
rect 6237 4123 6253 4187
rect 6317 4123 6333 4187
rect 6397 4123 6416 4187
rect 5416 4068 6416 4123
rect 5416 4004 5427 4068
rect 5491 4004 5507 4068
rect 5571 4004 5587 4068
rect 5651 4004 5667 4068
rect 5731 4004 6093 4068
rect 6157 4004 6173 4068
rect 6237 4004 6253 4068
rect 6317 4004 6333 4068
rect 6397 4004 6416 4068
rect 5416 -2464 6416 4004
rect 12130 16034 13130 22592
rect 12130 15970 12141 16034
rect 12205 15970 12221 16034
rect 12285 15970 12301 16034
rect 12365 15970 12381 16034
rect 12445 15970 12807 16034
rect 12871 15970 12887 16034
rect 12951 15970 12967 16034
rect 13031 15970 13047 16034
rect 13111 15970 13130 16034
rect 12130 15915 13130 15970
rect 12130 15851 12141 15915
rect 12205 15851 12221 15915
rect 12285 15851 12301 15915
rect 12365 15851 12381 15915
rect 12445 15851 12807 15915
rect 12871 15851 12887 15915
rect 12951 15851 12967 15915
rect 13031 15851 13047 15915
rect 13111 15851 13130 15915
rect 12130 4194 13130 15851
rect 12130 4130 12141 4194
rect 12205 4130 12221 4194
rect 12285 4130 12301 4194
rect 12365 4130 12381 4194
rect 12445 4130 12807 4194
rect 12871 4130 12887 4194
rect 12951 4130 12967 4194
rect 13031 4130 13047 4194
rect 13111 4130 13130 4194
rect 12130 4075 13130 4130
rect 12130 4011 12141 4075
rect 12205 4011 12221 4075
rect 12285 4011 12301 4075
rect 12365 4011 12381 4075
rect 12445 4011 12807 4075
rect 12871 4011 12887 4075
rect 12951 4011 12967 4075
rect 13031 4011 13047 4075
rect 13111 4011 13130 4075
rect 12130 -2464 13130 4011
use sky130_ef_ip__rc_osc_500k  sky130_ef_ip__rc_osc_500k_0
timestamp 1527949378
transform 0 -1 14561 1 0 4000
box 0 0 12242 10724
<< labels >>
flabel metal2 s 9006 20076 9118 21516 0 FreeSans 560 90 0 0 dout
port 1 nsew
flabel metal2 s 9650 20076 9762 21516 0 FreeSans 560 90 0 0 ena
port 2 nsew
flabel metal4 s 7440 16042 8197 23675 0 FreeSans 9600 90 0 0 vssd1
port 3 nsew
flabel metal4 s 10170 16042 10927 23675 0 FreeSans 9600 90 0 0 vccd1
port 4 nsew
flabel metal4 s 5416 -2464 6416 22592 0 FreeSans 9600 90 0 0 vdda1
port 5 nsew
flabel metal4 s 12130 -2464 13130 22592 0 FreeSans 9600 90 0 0 vssa1
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 18412 20556
<< end >>

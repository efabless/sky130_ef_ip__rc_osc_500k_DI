VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__rc_osc_500k_DI
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__rc_osc_500k_DI ;
  ORIGIN -18.585 -19.730 ;
  SIZE 54.360 BY 63.890 ;
  PIN dout
    ANTENNADIFFAREA 0.556800 ;
    PORT
      LAYER met2 ;
        RECT 45.030 82.095 45.590 89.295 ;
    END
  END dout
  PIN ena
    ANTENNAGATEAREA 0.858000 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 48.250 82.095 48.810 89.295 ;
    END
  END ena
  PIN vssd1
    ANTENNADIFFAREA 6.628900 ;
    PORT
      LAYER met4 ;
        RECT 37.200 80.210 40.985 118.375 ;
    END
  END vssd1
  PIN vccd1
    ANTENNADIFFAREA 4.280700 ;
    PORT
      LAYER met4 ;
        RECT 50.850 80.210 54.635 118.375 ;
    END
  END vccd1
  PIN vdda1
    ANTENNADIFFAREA 148.310989 ;
    PORT
      LAYER met4 ;
        RECT 27.080 -12.320 32.080 112.960 ;
    END
  END vdda1
  PIN vssa1
    ANTENNADIFFAREA 114.014595 ;
    PORT
      LAYER met4 ;
        RECT 60.650 -12.320 65.650 112.960 ;
    END
  END vssa1
  OBS
      LAYER nwell ;
        RECT 19.185 79.600 39.555 81.210 ;
        RECT 19.185 21.610 20.795 79.600 ;
        RECT 19.185 20.000 72.805 21.610 ;
      LAYER li1 ;
        RECT 19.625 20.430 72.340 80.755 ;
      LAYER met1 ;
        RECT 21.805 20.430 70.215 81.210 ;
      LAYER met2 ;
        RECT 24.325 81.815 44.750 83.295 ;
        RECT 45.870 81.815 47.970 83.295 ;
        RECT 49.090 81.815 67.465 83.295 ;
        RECT 24.325 20.000 67.465 81.815 ;
      LAYER met3 ;
        RECT 27.080 19.995 65.650 81.210 ;
      LAYER met4 ;
        RECT 44.815 31.555 54.955 57.335 ;
  END
END sky130_ef_ip__rc_osc_500k_DI
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__rc_osc_500k_DI
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__rc_osc_500k_DI ;
  ORIGIN 0.000 0.000 ;
  SIZE 92.060 BY 102.780 ;
  PIN dout
    ANTENNADIFFAREA 0.556800 ;
    PORT
      LAYER li1 ;
        RECT 45.840 79.525 46.880 79.695 ;
        RECT 48.410 79.105 48.950 79.275 ;
        RECT 41.855 71.530 42.315 71.700 ;
      LAYER mcon ;
        RECT 46.095 79.525 46.265 79.695 ;
        RECT 46.455 79.525 46.625 79.695 ;
        RECT 48.595 79.105 48.765 79.275 ;
        RECT 42.000 71.530 42.170 71.700 ;
      LAYER met1 ;
        RECT 43.895 79.675 47.375 79.880 ;
        RECT 43.895 79.550 45.155 79.675 ;
        RECT 43.895 79.435 44.740 79.550 ;
        RECT 45.860 79.495 46.860 79.675 ;
        RECT 47.170 79.140 47.375 79.675 ;
        RECT 48.430 79.140 48.930 79.305 ;
        RECT 47.170 79.075 48.930 79.140 ;
        RECT 47.170 78.935 48.875 79.075 ;
        RECT 41.875 71.535 42.295 71.730 ;
        RECT 41.865 71.305 43.135 71.535 ;
        RECT 41.865 71.270 43.225 71.305 ;
        RECT 42.865 70.325 43.225 71.270 ;
      LAYER via ;
        RECT 44.030 79.525 44.290 79.785 ;
        RECT 44.350 79.525 44.610 79.785 ;
        RECT 42.915 70.845 43.175 71.105 ;
        RECT 42.915 70.525 43.175 70.785 ;
      LAYER met2 ;
        RECT 45.030 101.050 45.590 107.580 ;
        RECT 44.320 100.910 45.590 101.050 ;
        RECT 44.320 81.210 44.460 100.910 ;
        RECT 45.030 100.380 45.590 100.910 ;
        RECT 43.655 80.210 44.655 81.210 ;
        RECT 44.010 79.830 44.230 80.210 ;
        RECT 43.845 79.485 44.790 79.830 ;
        RECT 44.010 77.870 44.230 79.485 ;
        RECT 42.940 77.650 44.230 77.870 ;
        RECT 42.940 71.255 43.160 77.650 ;
        RECT 42.815 70.375 43.275 71.255 ;
        RECT 42.940 70.370 43.160 70.375 ;
    END
  END dout
  PIN ena
    ANTENNAGATEAREA 0.858000 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 49.120 79.245 49.290 79.575 ;
        RECT 47.345 76.845 47.515 77.175 ;
        RECT 44.755 75.260 44.925 75.590 ;
        RECT 46.350 75.260 46.520 75.590 ;
        RECT 44.620 71.450 44.950 71.940 ;
        RECT 41.875 66.900 42.045 67.400 ;
        RECT 42.845 66.900 43.015 67.400 ;
        RECT 48.095 58.090 48.265 58.590 ;
        RECT 49.065 58.090 49.235 58.590 ;
      LAYER mcon ;
        RECT 49.120 79.325 49.290 79.495 ;
        RECT 47.345 76.925 47.515 77.095 ;
        RECT 44.755 75.340 44.925 75.510 ;
        RECT 46.350 75.340 46.520 75.510 ;
        RECT 44.700 71.610 44.870 71.780 ;
        RECT 41.875 67.065 42.045 67.235 ;
        RECT 42.845 67.065 43.015 67.235 ;
        RECT 48.095 58.255 48.265 58.425 ;
        RECT 49.065 58.255 49.235 58.425 ;
      LAYER met1 ;
        RECT 49.155 79.555 49.450 79.915 ;
        RECT 49.090 79.265 49.450 79.555 ;
        RECT 49.155 78.885 49.450 79.265 ;
        RECT 45.215 75.770 46.215 76.770 ;
        RECT 47.315 76.265 47.675 77.245 ;
        RECT 45.535 75.590 45.905 75.770 ;
        RECT 44.705 75.350 46.565 75.590 ;
        RECT 44.725 75.280 44.955 75.350 ;
        RECT 45.535 75.300 45.905 75.350 ;
        RECT 46.320 75.280 46.550 75.350 ;
        RECT 44.600 71.920 44.960 72.040 ;
        RECT 44.590 71.470 44.980 71.920 ;
        RECT 44.600 71.060 44.960 71.470 ;
        RECT 41.845 67.280 42.075 67.380 ;
        RECT 42.815 67.280 43.055 67.380 ;
        RECT 44.625 67.280 44.955 67.620 ;
        RECT 41.845 67.080 44.955 67.280 ;
        RECT 41.845 66.920 42.075 67.080 ;
        RECT 42.815 66.920 43.045 67.080 ;
        RECT 44.625 67.030 44.955 67.080 ;
        RECT 49.615 60.435 49.935 61.470 ;
        RECT 49.615 60.345 49.810 60.435 ;
        RECT 49.090 60.165 49.810 60.345 ;
        RECT 49.090 58.570 49.270 60.165 ;
        RECT 48.065 58.425 48.295 58.570 ;
        RECT 49.035 58.425 49.270 58.570 ;
        RECT 48.065 58.245 49.270 58.425 ;
        RECT 48.065 58.110 48.295 58.245 ;
        RECT 49.035 58.110 49.265 58.245 ;
      LAYER via ;
        RECT 49.175 79.590 49.435 79.850 ;
        RECT 49.175 79.270 49.435 79.530 ;
        RECT 49.175 78.950 49.435 79.210 ;
        RECT 47.365 76.785 47.625 77.045 ;
        RECT 47.365 76.465 47.625 76.725 ;
        RECT 45.590 75.420 45.850 75.680 ;
        RECT 44.650 71.580 44.910 71.840 ;
        RECT 44.650 71.260 44.910 71.520 ;
        RECT 44.660 67.195 44.920 67.455 ;
        RECT 49.645 61.140 49.905 61.400 ;
        RECT 49.645 60.820 49.905 61.080 ;
        RECT 49.645 60.500 49.905 60.760 ;
      LAYER met2 ;
        RECT 48.250 101.580 48.810 107.580 ;
        RECT 48.205 100.380 48.810 101.580 ;
        RECT 48.205 100.370 48.345 100.380 ;
        RECT 48.000 100.230 48.345 100.370 ;
        RECT 48.000 81.210 48.140 100.230 ;
        RECT 47.875 80.210 48.875 81.210 ;
        RECT 48.240 79.550 48.510 80.210 ;
        RECT 49.105 79.550 49.500 79.865 ;
        RECT 48.240 79.270 49.500 79.550 ;
        RECT 48.240 77.845 48.510 79.270 ;
        RECT 49.105 78.935 49.500 79.270 ;
        RECT 45.580 77.575 48.510 77.845 ;
        RECT 45.580 75.750 45.850 77.575 ;
        RECT 47.375 77.195 47.610 77.575 ;
        RECT 47.265 76.315 47.725 77.195 ;
        RECT 45.485 75.350 45.955 75.750 ;
        RECT 45.580 74.680 45.850 75.350 ;
        RECT 44.645 74.410 45.850 74.680 ;
        RECT 44.645 71.990 44.915 74.410 ;
        RECT 44.550 71.110 45.010 71.990 ;
        RECT 44.645 68.765 44.915 71.110 ;
        RECT 44.645 68.440 49.935 68.765 ;
        RECT 44.645 67.570 44.915 68.440 ;
        RECT 44.575 67.080 45.005 67.570 ;
        RECT 49.610 61.420 49.935 68.440 ;
        RECT 49.565 60.485 49.985 61.420 ;
        RECT 49.610 60.475 49.935 60.485 ;
    END
  END ena
  PIN vssd1
    ANTENNADIFFAREA 6.628900 ;
    PORT
      LAYER pwell ;
        RECT 41.920 78.370 44.110 80.380 ;
        RECT 47.740 78.405 49.930 80.415 ;
        RECT 41.245 74.320 41.975 75.650 ;
        RECT 42.875 74.420 45.565 76.430 ;
        RECT 41.185 70.830 43.295 72.840 ;
        RECT 43.920 70.830 45.650 72.560 ;
      LAYER li1 ;
        RECT 47.870 80.270 49.800 80.285 ;
        RECT 42.050 80.245 43.980 80.250 ;
        RECT 41.545 80.080 44.195 80.245 ;
        RECT 41.545 78.670 42.220 80.080 ;
        RECT 42.590 79.070 43.130 79.240 ;
        RECT 43.810 78.670 44.195 80.080 ;
        RECT 41.545 77.980 44.195 78.670 ;
        RECT 47.735 80.115 50.315 80.270 ;
        RECT 47.735 78.705 48.110 80.115 ;
        RECT 49.620 78.705 50.315 80.115 ;
        RECT 47.735 78.120 50.315 78.705 ;
        RECT 41.555 77.965 44.195 77.980 ;
        RECT 41.555 77.955 43.970 77.965 ;
        RECT 49.390 77.950 50.315 78.120 ;
        RECT 42.685 76.300 43.195 76.330 ;
        RECT 42.685 76.130 45.435 76.300 ;
        RECT 42.685 75.840 43.195 76.130 ;
        RECT 41.375 74.720 43.195 75.840 ;
        RECT 43.545 75.560 44.585 75.730 ;
        RECT 45.265 74.720 45.435 76.130 ;
        RECT 39.940 74.620 40.585 74.645 ;
        RECT 41.375 74.620 45.435 74.720 ;
        RECT 39.905 74.340 45.435 74.620 ;
        RECT 39.905 74.065 45.425 74.340 ;
        RECT 39.905 72.595 46.635 74.065 ;
        RECT 41.315 72.540 46.635 72.595 ;
        RECT 41.315 71.130 41.485 72.540 ;
        RECT 42.995 72.260 46.635 72.540 ;
        RECT 41.855 71.970 42.315 72.140 ;
        RECT 42.995 71.130 44.220 72.260 ;
        RECT 45.350 71.130 46.635 72.260 ;
        RECT 49.380 72.115 50.315 77.950 ;
        RECT 41.315 70.965 46.635 71.130 ;
        RECT 49.370 71.085 50.315 72.115 ;
        RECT 41.315 70.960 43.165 70.965 ;
        RECT 44.050 70.960 46.635 70.965 ;
        RECT 45.350 70.940 46.635 70.960 ;
      LAYER mcon ;
        RECT 42.775 79.070 42.945 79.240 ;
        RECT 41.615 78.180 42.145 79.070 ;
        RECT 42.765 78.440 42.935 78.610 ;
        RECT 42.765 78.080 42.935 78.250 ;
        RECT 43.800 75.560 43.970 75.730 ;
        RECT 44.160 75.560 44.330 75.730 ;
        RECT 42.185 75.000 42.715 75.530 ;
        RECT 40.000 73.280 40.530 74.530 ;
        RECT 42.000 71.970 42.170 72.140 ;
        RECT 45.555 71.320 46.445 71.850 ;
        RECT 49.575 71.330 50.105 71.860 ;
      LAYER met1 ;
        RECT 37.200 79.320 40.985 81.210 ;
        RECT 39.985 79.195 40.985 79.320 ;
        RECT 39.985 78.145 42.225 79.195 ;
        RECT 42.610 79.040 43.110 79.270 ;
        RECT 42.610 78.145 43.080 79.040 ;
        RECT 39.985 76.710 43.080 78.145 ;
        RECT 39.985 76.640 43.090 76.710 ;
        RECT 39.985 75.980 43.105 76.640 ;
        RECT 39.985 75.750 44.575 75.980 ;
        RECT 39.985 75.740 43.165 75.750 ;
        RECT 39.985 75.710 43.105 75.740 ;
        RECT 39.910 73.105 40.615 74.705 ;
        RECT 42.105 74.400 43.105 75.710 ;
        RECT 43.565 75.530 44.565 75.750 ;
        RECT 40.030 72.265 40.390 72.315 ;
        RECT 40.030 71.955 42.295 72.265 ;
        RECT 40.030 71.335 40.390 71.955 ;
        RECT 41.875 71.940 42.295 71.955 ;
        RECT 45.340 71.085 50.305 72.115 ;
      LAYER via ;
        RECT 37.260 80.915 37.520 81.175 ;
        RECT 37.580 80.915 37.840 81.175 ;
        RECT 37.900 80.915 38.160 81.175 ;
        RECT 38.220 80.915 38.480 81.175 ;
        RECT 39.100 80.915 39.360 81.175 ;
        RECT 39.420 80.915 39.680 81.175 ;
        RECT 39.740 80.915 40.000 81.175 ;
        RECT 40.630 80.910 40.890 81.170 ;
        RECT 37.260 80.465 37.520 80.725 ;
        RECT 37.580 80.465 37.840 80.725 ;
        RECT 37.900 80.465 38.160 80.725 ;
        RECT 38.220 80.465 38.480 80.725 ;
        RECT 39.100 80.465 39.360 80.725 ;
        RECT 39.420 80.465 39.680 80.725 ;
        RECT 39.740 80.465 40.000 80.725 ;
        RECT 40.630 80.460 40.890 80.720 ;
        RECT 40.155 77.175 40.415 77.435 ;
        RECT 40.155 76.855 40.415 77.115 ;
        RECT 40.155 76.535 40.415 76.795 ;
        RECT 40.155 76.215 40.415 76.475 ;
        RECT 40.155 75.895 40.415 76.155 ;
        RECT 39.975 73.295 40.555 74.515 ;
        RECT 40.080 71.855 40.340 72.115 ;
        RECT 40.080 71.535 40.340 71.795 ;
      LAYER met2 ;
        RECT 37.200 80.210 40.985 81.210 ;
        RECT 39.935 74.645 40.595 77.590 ;
        RECT 39.890 73.165 40.635 74.645 ;
        RECT 39.935 71.315 40.595 73.165 ;
      LAYER via2 ;
        RECT 37.275 80.885 37.555 81.165 ;
        RECT 37.675 80.885 37.955 81.165 ;
        RECT 38.075 80.885 38.355 81.165 ;
        RECT 38.475 80.885 38.755 81.165 ;
        RECT 39.105 80.885 39.385 81.165 ;
        RECT 39.505 80.885 39.785 81.165 ;
        RECT 39.905 80.885 40.185 81.165 ;
        RECT 40.305 80.885 40.585 81.165 ;
        RECT 37.275 80.290 37.555 80.570 ;
        RECT 37.675 80.290 37.955 80.570 ;
        RECT 38.075 80.290 38.355 80.570 ;
        RECT 38.475 80.290 38.755 80.570 ;
        RECT 39.105 80.290 39.385 80.570 ;
        RECT 39.505 80.290 39.785 80.570 ;
        RECT 39.905 80.290 40.185 80.570 ;
        RECT 40.305 80.290 40.585 80.570 ;
      LAYER met3 ;
        RECT 37.200 80.210 40.985 81.210 ;
      LAYER via3 ;
        RECT 37.255 80.865 37.575 81.185 ;
        RECT 37.655 80.865 37.975 81.185 ;
        RECT 38.055 80.865 38.375 81.185 ;
        RECT 38.455 80.865 38.775 81.185 ;
        RECT 39.085 80.865 39.405 81.185 ;
        RECT 39.485 80.865 39.805 81.185 ;
        RECT 39.885 80.865 40.205 81.185 ;
        RECT 40.285 80.865 40.605 81.185 ;
        RECT 37.255 80.270 37.575 80.590 ;
        RECT 37.655 80.270 37.975 80.590 ;
        RECT 38.055 80.270 38.375 80.590 ;
        RECT 38.455 80.270 38.775 80.590 ;
        RECT 39.085 80.270 39.405 80.590 ;
        RECT 39.485 80.270 39.805 80.590 ;
        RECT 39.885 80.270 40.205 80.590 ;
        RECT 40.285 80.270 40.605 80.590 ;
      LAYER met4 ;
        RECT 37.200 80.210 40.985 118.375 ;
    END
  END vssd1
  PIN vccd1
    ANTENNADIFFAREA 4.280700 ;
    PORT
      LAYER nwell ;
        RECT 44.760 78.335 47.600 80.445 ;
        RECT 45.840 78.065 47.600 78.335 ;
        RECT 45.950 76.480 48.210 78.065 ;
        RECT 45.655 74.370 48.495 76.480 ;
      LAYER li1 ;
        RECT 47.150 80.265 47.525 80.270 ;
        RECT 44.940 80.245 47.525 80.265 ;
        RECT 44.730 80.095 47.525 80.245 ;
        RECT 44.730 78.690 45.110 80.095 ;
        RECT 45.840 79.085 46.880 79.255 ;
        RECT 47.150 78.690 47.525 80.095 ;
        RECT 44.730 77.975 47.525 78.690 ;
        RECT 44.730 77.965 45.105 77.975 ;
        RECT 45.825 77.885 47.525 77.975 ;
        RECT 45.825 77.860 48.675 77.885 ;
        RECT 46.130 77.715 48.675 77.860 ;
        RECT 46.130 76.305 46.300 77.715 ;
        RECT 46.670 77.145 47.130 77.315 ;
        RECT 47.860 76.305 48.675 77.715 ;
        RECT 46.130 76.300 48.675 76.305 ;
        RECT 45.835 76.130 48.675 76.300 ;
        RECT 45.835 74.720 46.005 76.130 ;
        RECT 48.145 75.850 48.675 76.130 ;
        RECT 46.735 75.560 47.775 75.730 ;
        RECT 48.145 75.060 49.135 75.850 ;
        RECT 48.145 74.720 48.675 75.060 ;
        RECT 45.835 74.330 48.675 74.720 ;
        RECT 44.100 57.920 44.560 58.090 ;
      LAYER mcon ;
        RECT 46.095 79.085 46.265 79.255 ;
        RECT 46.455 79.085 46.625 79.255 ;
        RECT 45.910 78.075 46.800 78.605 ;
        RECT 46.815 77.145 46.985 77.315 ;
        RECT 46.990 75.560 47.160 75.730 ;
        RECT 47.350 75.560 47.520 75.730 ;
        RECT 48.465 75.170 48.995 75.700 ;
        RECT 44.245 57.920 44.415 58.090 ;
      LAYER met1 ;
        RECT 50.850 79.320 54.635 81.210 ;
        RECT 45.860 79.055 46.860 79.285 ;
        RECT 45.865 78.705 46.855 79.055 ;
        RECT 45.805 78.575 46.905 78.705 ;
        RECT 50.850 78.575 51.850 79.320 ;
        RECT 45.805 77.975 51.850 78.575 ;
        RECT 45.865 77.515 51.850 77.975 ;
        RECT 46.695 77.345 47.105 77.515 ;
        RECT 46.690 77.115 47.110 77.345 ;
        RECT 48.135 75.930 51.850 77.515 ;
        RECT 46.755 75.775 51.850 75.930 ;
        RECT 46.755 75.700 49.135 75.775 ;
        RECT 46.755 75.530 47.755 75.700 ;
        RECT 41.425 74.030 41.920 75.090 ;
        RECT 48.135 74.030 49.135 75.700 ;
        RECT 41.425 73.220 49.135 74.030 ;
        RECT 41.425 73.190 41.920 73.220 ;
        RECT 41.445 57.975 41.940 59.410 ;
        RECT 44.120 57.975 44.540 58.120 ;
        RECT 41.445 57.890 44.540 57.975 ;
        RECT 41.445 57.555 44.475 57.890 ;
        RECT 41.445 57.510 41.940 57.555 ;
      LAYER via ;
        RECT 50.930 80.915 51.190 81.175 ;
        RECT 51.250 80.915 51.510 81.175 ;
        RECT 51.570 80.915 51.830 81.175 ;
        RECT 51.890 80.915 52.150 81.175 ;
        RECT 52.770 80.915 53.030 81.175 ;
        RECT 53.090 80.915 53.350 81.175 ;
        RECT 53.410 80.915 53.670 81.175 ;
        RECT 54.300 80.910 54.560 81.170 ;
        RECT 50.930 80.465 51.190 80.725 ;
        RECT 51.250 80.465 51.510 80.725 ;
        RECT 51.570 80.465 51.830 80.725 ;
        RECT 51.890 80.465 52.150 80.725 ;
        RECT 52.770 80.465 53.030 80.725 ;
        RECT 53.090 80.465 53.350 80.725 ;
        RECT 53.410 80.465 53.670 80.725 ;
        RECT 54.300 80.460 54.560 80.720 ;
        RECT 41.545 74.650 41.805 74.910 ;
        RECT 41.545 74.330 41.805 74.590 ;
        RECT 41.545 74.010 41.805 74.270 ;
        RECT 41.545 73.690 41.805 73.950 ;
        RECT 41.545 73.370 41.805 73.630 ;
        RECT 41.565 58.970 41.825 59.230 ;
        RECT 41.565 58.650 41.825 58.910 ;
        RECT 41.565 58.330 41.825 58.590 ;
        RECT 41.565 58.010 41.825 58.270 ;
        RECT 41.565 57.690 41.825 57.950 ;
      LAYER met2 ;
        RECT 50.850 80.210 54.635 81.210 ;
        RECT 41.375 73.240 41.970 75.040 ;
        RECT 41.435 59.360 41.925 73.240 ;
        RECT 41.395 57.560 41.990 59.360 ;
      LAYER via2 ;
        RECT 50.925 80.885 51.205 81.165 ;
        RECT 51.325 80.885 51.605 81.165 ;
        RECT 51.725 80.885 52.005 81.165 ;
        RECT 52.125 80.885 52.405 81.165 ;
        RECT 52.755 80.885 53.035 81.165 ;
        RECT 53.155 80.885 53.435 81.165 ;
        RECT 53.555 80.885 53.835 81.165 ;
        RECT 53.955 80.885 54.235 81.165 ;
        RECT 50.925 80.290 51.205 80.570 ;
        RECT 51.325 80.290 51.605 80.570 ;
        RECT 51.725 80.290 52.005 80.570 ;
        RECT 52.125 80.290 52.405 80.570 ;
        RECT 52.755 80.290 53.035 80.570 ;
        RECT 53.155 80.290 53.435 80.570 ;
        RECT 53.555 80.290 53.835 80.570 ;
        RECT 53.955 80.290 54.235 80.570 ;
      LAYER met3 ;
        RECT 50.850 80.210 54.635 81.210 ;
      LAYER via3 ;
        RECT 50.905 80.865 51.225 81.185 ;
        RECT 51.305 80.865 51.625 81.185 ;
        RECT 51.705 80.865 52.025 81.185 ;
        RECT 52.105 80.865 52.425 81.185 ;
        RECT 52.735 80.865 53.055 81.185 ;
        RECT 53.135 80.865 53.455 81.185 ;
        RECT 53.535 80.865 53.855 81.185 ;
        RECT 53.935 80.865 54.255 81.185 ;
        RECT 50.905 80.270 51.225 80.590 ;
        RECT 51.305 80.270 51.625 80.590 ;
        RECT 51.705 80.270 52.025 80.590 ;
        RECT 52.105 80.270 52.425 80.590 ;
        RECT 52.735 80.270 53.055 80.590 ;
        RECT 53.135 80.270 53.455 80.590 ;
        RECT 53.535 80.270 53.855 80.590 ;
        RECT 53.935 80.270 54.255 80.590 ;
      LAYER met4 ;
        RECT 50.850 80.210 54.635 118.375 ;
    END
  END vccd1
  PIN vdda1
    ANTENNADIFFAREA 148.310989 ;
    PORT
      LAYER nwell ;
        RECT 19.185 79.600 39.555 81.210 ;
        RECT 19.185 21.610 20.795 79.600 ;
        RECT 37.945 70.450 39.555 79.600 ;
        RECT 52.455 79.600 72.805 81.210 ;
        RECT 52.455 70.450 54.065 79.600 ;
        RECT 37.945 68.840 54.065 70.450 ;
        RECT 44.265 65.650 52.115 68.840 ;
        RECT 44.255 62.570 52.115 65.650 ;
        RECT 39.240 55.590 46.025 59.940 ;
        RECT 39.245 30.950 46.025 55.590 ;
        RECT 71.195 21.610 72.805 79.600 ;
        RECT 19.185 20.000 72.805 21.610 ;
      LAYER li1 ;
        RECT 19.625 80.745 20.340 80.755 ;
        RECT 19.625 80.230 39.150 80.745 ;
        RECT 19.625 21.050 20.340 80.230 ;
        RECT 38.340 70.020 39.150 80.230 ;
        RECT 52.720 80.230 72.340 80.745 ;
        RECT 52.720 70.020 53.340 80.230 ;
        RECT 38.340 69.275 53.340 70.020 ;
        RECT 44.295 68.150 51.045 68.780 ;
        RECT 44.295 68.140 48.165 68.150 ;
        RECT 44.295 66.180 44.835 68.140 ;
        RECT 47.095 66.210 48.165 68.140 ;
        RECT 49.070 66.710 49.530 66.880 ;
        RECT 50.425 66.210 51.045 68.150 ;
        RECT 47.095 66.180 51.045 66.210 ;
        RECT 44.295 65.090 51.045 66.180 ;
        RECT 44.295 63.170 44.835 65.090 ;
        RECT 47.085 63.170 48.165 65.090 ;
        RECT 49.070 64.420 49.530 64.590 ;
        RECT 50.425 63.170 51.045 65.090 ;
        RECT 44.295 62.540 51.045 63.170 ;
        RECT 51.525 61.560 53.190 68.580 ;
        RECT 42.050 59.500 46.250 60.045 ;
        RECT 42.050 59.425 46.255 59.500 ;
        RECT 39.045 59.380 46.255 59.425 ;
        RECT 39.045 57.825 43.195 59.380 ;
        RECT 39.045 55.200 39.840 57.825 ;
        RECT 42.055 57.420 43.195 57.825 ;
        RECT 45.460 57.420 46.255 59.380 ;
        RECT 42.055 57.250 46.255 57.420 ;
        RECT 42.055 55.445 43.185 57.250 ;
        RECT 42.050 55.200 43.185 55.445 ;
        RECT 45.460 55.200 46.255 57.250 ;
        RECT 39.045 55.030 46.255 55.200 ;
        RECT 39.045 53.070 39.840 55.030 ;
        RECT 40.710 54.360 41.170 54.530 ;
        RECT 42.050 54.075 43.195 55.030 ;
        RECT 42.055 53.070 43.195 54.075 ;
        RECT 45.460 53.070 46.255 55.030 ;
        RECT 39.045 52.900 46.255 53.070 ;
        RECT 39.045 52.120 39.840 52.900 ;
        RECT 42.055 52.365 43.185 52.900 ;
        RECT 42.050 52.120 43.185 52.365 ;
        RECT 45.460 52.120 46.255 52.900 ;
        RECT 39.045 51.950 46.255 52.120 ;
        RECT 39.045 49.990 39.840 51.950 ;
        RECT 40.710 51.280 41.170 51.450 ;
        RECT 42.050 50.995 43.195 51.950 ;
        RECT 42.055 49.990 43.195 50.995 ;
        RECT 45.460 49.990 46.255 51.950 ;
        RECT 39.045 49.820 46.255 49.990 ;
        RECT 39.045 49.040 39.840 49.820 ;
        RECT 42.055 49.285 43.185 49.820 ;
        RECT 42.050 49.040 43.185 49.285 ;
        RECT 45.460 49.040 46.255 49.820 ;
        RECT 39.045 48.870 46.255 49.040 ;
        RECT 39.045 46.910 39.840 48.870 ;
        RECT 40.710 48.200 41.170 48.370 ;
        RECT 42.050 47.915 43.195 48.870 ;
        RECT 42.055 46.910 43.195 47.915 ;
        RECT 45.460 46.910 46.255 48.870 ;
        RECT 39.045 46.740 46.255 46.910 ;
        RECT 39.045 45.960 39.840 46.740 ;
        RECT 42.055 46.205 43.185 46.740 ;
        RECT 42.050 45.960 43.185 46.205 ;
        RECT 45.460 45.960 46.255 46.740 ;
        RECT 39.045 45.790 46.255 45.960 ;
        RECT 39.045 43.830 39.840 45.790 ;
        RECT 40.710 45.120 41.170 45.290 ;
        RECT 42.050 44.835 43.195 45.790 ;
        RECT 42.055 43.830 43.195 44.835 ;
        RECT 45.460 43.830 46.255 45.790 ;
        RECT 39.045 43.660 46.255 43.830 ;
        RECT 39.045 42.880 39.840 43.660 ;
        RECT 42.055 43.125 43.185 43.660 ;
        RECT 42.050 42.880 43.185 43.125 ;
        RECT 45.460 42.880 46.255 43.660 ;
        RECT 39.045 42.710 46.255 42.880 ;
        RECT 39.045 40.750 39.840 42.710 ;
        RECT 40.710 42.040 41.170 42.210 ;
        RECT 42.050 41.755 43.195 42.710 ;
        RECT 42.055 40.750 43.195 41.755 ;
        RECT 45.460 40.750 46.255 42.710 ;
        RECT 39.045 40.580 46.255 40.750 ;
        RECT 39.045 39.800 39.840 40.580 ;
        RECT 42.055 40.045 43.185 40.580 ;
        RECT 42.050 39.800 43.185 40.045 ;
        RECT 45.460 39.800 46.255 40.580 ;
        RECT 39.045 39.630 46.255 39.800 ;
        RECT 39.045 37.670 39.840 39.630 ;
        RECT 40.710 38.960 41.170 39.130 ;
        RECT 42.050 38.675 43.195 39.630 ;
        RECT 42.055 37.670 43.195 38.675 ;
        RECT 45.460 37.670 46.255 39.630 ;
        RECT 39.045 37.500 46.255 37.670 ;
        RECT 39.045 36.720 39.840 37.500 ;
        RECT 42.055 36.965 43.185 37.500 ;
        RECT 42.050 36.720 43.185 36.965 ;
        RECT 45.460 36.720 46.255 37.500 ;
        RECT 39.045 36.550 46.255 36.720 ;
        RECT 39.045 34.590 39.840 36.550 ;
        RECT 40.710 35.880 41.170 36.050 ;
        RECT 42.050 35.595 43.195 36.550 ;
        RECT 42.055 34.590 43.195 35.595 ;
        RECT 45.460 34.590 46.255 36.550 ;
        RECT 39.045 34.420 46.255 34.590 ;
        RECT 39.045 33.640 39.840 34.420 ;
        RECT 42.055 33.885 43.185 34.420 ;
        RECT 42.050 33.640 43.185 33.885 ;
        RECT 45.460 33.640 46.255 34.420 ;
        RECT 39.045 33.470 46.255 33.640 ;
        RECT 39.045 31.510 39.840 33.470 ;
        RECT 40.710 32.800 41.170 32.970 ;
        RECT 42.050 32.515 43.195 33.470 ;
        RECT 44.100 32.800 44.560 32.970 ;
        RECT 42.055 31.510 43.195 32.515 ;
        RECT 45.460 31.510 46.255 33.470 ;
        RECT 39.045 30.905 46.255 31.510 ;
        RECT 39.050 30.670 46.245 30.905 ;
        RECT 55.055 22.670 57.215 23.020 ;
        RECT 71.810 21.050 72.340 80.230 ;
        RECT 19.625 20.430 72.340 21.050 ;
      LAYER mcon ;
        RECT 24.545 80.405 24.715 80.575 ;
        RECT 24.905 80.405 25.075 80.575 ;
        RECT 25.265 80.405 25.435 80.575 ;
        RECT 25.625 80.405 25.795 80.575 ;
        RECT 25.985 80.405 26.155 80.575 ;
        RECT 26.345 80.405 26.515 80.575 ;
        RECT 26.705 80.405 26.875 80.575 ;
        RECT 27.065 80.405 27.235 80.575 ;
        RECT 27.425 80.405 27.595 80.575 ;
        RECT 27.785 80.405 27.955 80.575 ;
        RECT 28.145 80.405 28.315 80.575 ;
        RECT 28.505 80.405 28.675 80.575 ;
        RECT 28.865 80.405 29.035 80.575 ;
        RECT 29.225 80.405 29.395 80.575 ;
        RECT 29.585 80.405 29.755 80.575 ;
        RECT 29.945 80.405 30.115 80.575 ;
        RECT 30.305 80.405 30.475 80.575 ;
        RECT 30.665 80.405 30.835 80.575 ;
        RECT 31.025 80.405 31.195 80.575 ;
        RECT 31.385 80.405 31.555 80.575 ;
        RECT 31.745 80.405 31.915 80.575 ;
        RECT 32.105 80.405 32.275 80.575 ;
        RECT 32.465 80.405 32.635 80.575 ;
        RECT 32.825 80.405 32.995 80.575 ;
        RECT 33.185 80.405 33.355 80.575 ;
        RECT 33.545 80.405 33.715 80.575 ;
        RECT 33.905 80.405 34.075 80.575 ;
        RECT 38.555 77.055 38.725 77.225 ;
        RECT 38.555 76.695 38.725 76.865 ;
        RECT 38.555 76.335 38.725 76.505 ;
        RECT 38.555 75.975 38.725 76.145 ;
        RECT 38.555 75.615 38.725 75.785 ;
        RECT 38.555 75.255 38.725 75.425 ;
        RECT 38.555 74.895 38.725 75.065 ;
        RECT 38.555 74.535 38.725 74.705 ;
        RECT 38.555 74.175 38.725 74.345 ;
        RECT 38.555 73.815 38.725 73.985 ;
        RECT 38.555 73.455 38.725 73.625 ;
        RECT 38.555 73.095 38.725 73.265 ;
        RECT 38.555 72.735 38.725 72.905 ;
        RECT 38.555 72.375 38.725 72.545 ;
        RECT 38.555 72.015 38.725 72.185 ;
        RECT 38.555 71.655 38.725 71.825 ;
        RECT 38.555 71.295 38.725 71.465 ;
        RECT 38.555 70.935 38.725 71.105 ;
        RECT 38.555 70.575 38.725 70.745 ;
        RECT 38.555 70.215 38.725 70.385 ;
        RECT 38.740 69.475 38.910 69.645 ;
        RECT 39.100 69.475 39.270 69.645 ;
        RECT 39.460 69.475 39.630 69.645 ;
        RECT 39.820 69.475 39.990 69.645 ;
        RECT 40.180 69.475 40.350 69.645 ;
        RECT 40.540 69.475 40.710 69.645 ;
        RECT 40.900 69.475 41.070 69.645 ;
        RECT 41.260 69.475 41.430 69.645 ;
        RECT 41.620 69.475 41.790 69.645 ;
        RECT 41.980 69.475 42.150 69.645 ;
        RECT 42.340 69.475 42.510 69.645 ;
        RECT 42.700 69.475 42.870 69.645 ;
        RECT 43.060 69.475 43.230 69.645 ;
        RECT 43.420 69.475 43.590 69.645 ;
        RECT 43.780 69.475 43.950 69.645 ;
        RECT 44.140 69.475 44.310 69.645 ;
        RECT 44.500 69.475 44.670 69.645 ;
        RECT 44.860 69.475 45.030 69.645 ;
        RECT 45.220 69.475 45.390 69.645 ;
        RECT 45.580 69.475 45.750 69.645 ;
        RECT 45.940 69.475 46.110 69.645 ;
        RECT 46.300 69.475 46.470 69.645 ;
        RECT 46.660 69.475 46.830 69.645 ;
        RECT 47.020 69.475 47.190 69.645 ;
        RECT 47.380 69.475 47.550 69.645 ;
        RECT 47.740 69.475 47.910 69.645 ;
        RECT 48.100 69.475 48.270 69.645 ;
        RECT 48.460 69.475 48.630 69.645 ;
        RECT 48.820 69.475 48.990 69.645 ;
        RECT 49.180 69.475 49.350 69.645 ;
        RECT 49.540 69.475 49.710 69.645 ;
        RECT 49.900 69.475 50.070 69.645 ;
        RECT 50.260 69.475 50.430 69.645 ;
        RECT 50.620 69.475 50.790 69.645 ;
        RECT 50.980 69.475 51.150 69.645 ;
        RECT 51.340 69.475 51.510 69.645 ;
        RECT 51.700 69.475 51.870 69.645 ;
        RECT 52.060 69.475 52.230 69.645 ;
        RECT 52.420 69.475 52.590 69.645 ;
        RECT 52.780 69.475 52.950 69.645 ;
        RECT 49.990 68.390 50.160 68.560 ;
        RECT 50.350 68.390 50.520 68.560 ;
        RECT 50.710 68.390 50.880 68.560 ;
        RECT 49.215 66.710 49.385 66.880 ;
        RECT 49.265 65.395 50.875 65.925 ;
        RECT 49.215 64.420 49.385 64.590 ;
        RECT 49.935 62.760 50.105 62.930 ;
        RECT 50.295 62.760 50.465 62.930 ;
        RECT 50.655 62.760 50.825 62.930 ;
        RECT 51.555 61.565 53.165 68.575 ;
        RECT 39.240 58.975 39.410 59.145 ;
        RECT 39.240 58.615 39.410 58.785 ;
        RECT 39.240 58.255 39.410 58.425 ;
        RECT 39.240 57.895 39.410 58.065 ;
        RECT 39.240 57.535 39.410 57.705 ;
        RECT 39.240 57.175 39.410 57.345 ;
        RECT 39.240 56.815 39.410 56.985 ;
        RECT 39.240 56.455 39.410 56.625 ;
        RECT 39.240 56.095 39.410 56.265 ;
        RECT 39.240 55.735 39.410 55.905 ;
        RECT 39.240 55.375 39.410 55.545 ;
        RECT 39.240 55.015 39.410 55.185 ;
        RECT 39.240 54.655 39.410 54.825 ;
        RECT 39.240 54.295 39.410 54.465 ;
        RECT 40.855 54.360 41.025 54.530 ;
        RECT 39.240 53.935 39.410 54.105 ;
        RECT 42.175 54.135 43.065 55.385 ;
        RECT 39.240 53.575 39.410 53.745 ;
        RECT 39.240 53.215 39.410 53.385 ;
        RECT 39.240 52.855 39.410 53.025 ;
        RECT 39.240 52.495 39.410 52.665 ;
        RECT 39.240 52.135 39.410 52.305 ;
        RECT 39.240 51.775 39.410 51.945 ;
        RECT 39.240 51.415 39.410 51.585 ;
        RECT 40.855 51.280 41.025 51.450 ;
        RECT 39.240 51.055 39.410 51.225 ;
        RECT 42.175 51.055 43.065 52.305 ;
        RECT 39.240 50.695 39.410 50.865 ;
        RECT 39.240 50.335 39.410 50.505 ;
        RECT 39.240 49.975 39.410 50.145 ;
        RECT 39.240 49.615 39.410 49.785 ;
        RECT 39.240 49.255 39.410 49.425 ;
        RECT 39.240 48.895 39.410 49.065 ;
        RECT 39.240 48.535 39.410 48.705 ;
        RECT 39.240 48.175 39.410 48.345 ;
        RECT 40.855 48.200 41.025 48.370 ;
        RECT 39.240 47.815 39.410 47.985 ;
        RECT 42.175 47.975 43.065 49.225 ;
        RECT 39.240 47.455 39.410 47.625 ;
        RECT 39.240 47.095 39.410 47.265 ;
        RECT 39.240 46.735 39.410 46.905 ;
        RECT 39.240 46.375 39.410 46.545 ;
        RECT 39.240 46.015 39.410 46.185 ;
        RECT 39.240 45.655 39.410 45.825 ;
        RECT 39.240 45.295 39.410 45.465 ;
        RECT 40.855 45.120 41.025 45.290 ;
        RECT 39.240 44.935 39.410 45.105 ;
        RECT 42.175 44.895 43.065 46.145 ;
        RECT 39.240 44.575 39.410 44.745 ;
        RECT 39.240 44.215 39.410 44.385 ;
        RECT 39.240 43.855 39.410 44.025 ;
        RECT 39.240 43.495 39.410 43.665 ;
        RECT 39.240 43.135 39.410 43.305 ;
        RECT 39.240 42.775 39.410 42.945 ;
        RECT 39.240 42.415 39.410 42.585 ;
        RECT 39.240 42.055 39.410 42.225 ;
        RECT 40.855 42.040 41.025 42.210 ;
        RECT 39.240 41.695 39.410 41.865 ;
        RECT 42.175 41.815 43.065 43.065 ;
        RECT 39.240 41.335 39.410 41.505 ;
        RECT 39.240 40.975 39.410 41.145 ;
        RECT 39.240 40.615 39.410 40.785 ;
        RECT 39.240 40.255 39.410 40.425 ;
        RECT 39.240 39.895 39.410 40.065 ;
        RECT 39.240 39.535 39.410 39.705 ;
        RECT 39.240 39.175 39.410 39.345 ;
        RECT 39.240 38.815 39.410 38.985 ;
        RECT 40.855 38.960 41.025 39.130 ;
        RECT 42.175 38.735 43.065 39.985 ;
        RECT 39.240 38.455 39.410 38.625 ;
        RECT 39.240 38.095 39.410 38.265 ;
        RECT 39.240 37.735 39.410 37.905 ;
        RECT 39.240 37.375 39.410 37.545 ;
        RECT 39.240 37.015 39.410 37.185 ;
        RECT 39.240 36.655 39.410 36.825 ;
        RECT 39.240 36.295 39.410 36.465 ;
        RECT 39.240 35.935 39.410 36.105 ;
        RECT 40.855 35.880 41.025 36.050 ;
        RECT 39.240 35.575 39.410 35.745 ;
        RECT 42.175 35.655 43.065 36.905 ;
        RECT 39.240 35.215 39.410 35.385 ;
        RECT 39.240 34.855 39.410 35.025 ;
        RECT 39.240 34.495 39.410 34.665 ;
        RECT 39.240 34.135 39.410 34.305 ;
        RECT 39.240 33.775 39.410 33.945 ;
        RECT 39.240 33.415 39.410 33.585 ;
        RECT 39.240 33.055 39.410 33.225 ;
        RECT 39.240 32.695 39.410 32.865 ;
        RECT 40.855 32.800 41.025 32.970 ;
        RECT 42.175 32.575 43.065 33.825 ;
        RECT 44.245 32.800 44.415 32.970 ;
        RECT 39.240 32.335 39.410 32.505 ;
        RECT 39.240 31.975 39.410 32.145 ;
        RECT 39.240 31.615 39.410 31.785 ;
        RECT 39.240 31.255 39.410 31.425 ;
        RECT 55.155 22.760 55.325 22.930 ;
        RECT 55.515 22.760 55.685 22.930 ;
        RECT 55.875 22.760 56.045 22.930 ;
        RECT 56.235 22.760 56.405 22.930 ;
        RECT 56.595 22.760 56.765 22.930 ;
        RECT 56.955 22.760 57.125 22.930 ;
        RECT 34.500 20.675 34.670 20.845 ;
        RECT 34.860 20.675 35.030 20.845 ;
        RECT 35.220 20.675 35.390 20.845 ;
        RECT 35.580 20.675 35.750 20.845 ;
        RECT 35.940 20.675 36.110 20.845 ;
        RECT 36.300 20.675 36.470 20.845 ;
        RECT 36.660 20.675 36.830 20.845 ;
        RECT 37.020 20.675 37.190 20.845 ;
        RECT 37.380 20.675 37.550 20.845 ;
        RECT 37.740 20.675 37.910 20.845 ;
        RECT 38.100 20.675 38.270 20.845 ;
        RECT 38.460 20.675 38.630 20.845 ;
        RECT 38.820 20.675 38.990 20.845 ;
        RECT 39.180 20.675 39.350 20.845 ;
        RECT 39.540 20.675 39.710 20.845 ;
        RECT 39.900 20.675 40.070 20.845 ;
        RECT 40.260 20.675 40.430 20.845 ;
        RECT 40.620 20.675 40.790 20.845 ;
        RECT 40.980 20.675 41.150 20.845 ;
        RECT 41.340 20.675 41.510 20.845 ;
        RECT 41.700 20.675 41.870 20.845 ;
        RECT 42.060 20.675 42.230 20.845 ;
        RECT 42.420 20.675 42.590 20.845 ;
        RECT 42.780 20.675 42.950 20.845 ;
        RECT 43.140 20.675 43.310 20.845 ;
        RECT 43.500 20.675 43.670 20.845 ;
        RECT 43.860 20.675 44.030 20.845 ;
        RECT 44.220 20.675 44.390 20.845 ;
        RECT 44.580 20.675 44.750 20.845 ;
        RECT 44.940 20.675 45.110 20.845 ;
        RECT 45.300 20.675 45.470 20.845 ;
        RECT 45.660 20.675 45.830 20.845 ;
        RECT 46.020 20.675 46.190 20.845 ;
        RECT 46.380 20.675 46.550 20.845 ;
        RECT 46.740 20.675 46.910 20.845 ;
        RECT 47.100 20.675 47.270 20.845 ;
        RECT 47.460 20.675 47.630 20.845 ;
        RECT 47.820 20.675 47.990 20.845 ;
        RECT 48.180 20.675 48.350 20.845 ;
        RECT 48.540 20.675 48.710 20.845 ;
        RECT 48.900 20.675 49.070 20.845 ;
        RECT 49.260 20.675 49.430 20.845 ;
        RECT 49.620 20.675 49.790 20.845 ;
        RECT 49.980 20.675 50.150 20.845 ;
        RECT 50.340 20.675 50.510 20.845 ;
        RECT 50.700 20.675 50.870 20.845 ;
        RECT 51.060 20.675 51.230 20.845 ;
        RECT 51.420 20.675 51.590 20.845 ;
        RECT 51.780 20.675 51.950 20.845 ;
        RECT 52.140 20.675 52.310 20.845 ;
        RECT 52.500 20.675 52.670 20.845 ;
      LAYER met1 ;
        RECT 24.375 80.740 34.245 80.760 ;
        RECT 24.315 80.240 34.305 80.740 ;
        RECT 24.375 80.220 34.245 80.240 ;
        RECT 37.685 70.070 38.935 77.470 ;
        RECT 37.685 69.185 53.345 70.070 ;
        RECT 51.225 68.790 53.345 69.185 ;
        RECT 49.825 68.160 53.345 68.790 ;
        RECT 49.090 66.890 49.510 66.910 ;
        RECT 49.085 66.570 49.515 66.890 ;
        RECT 50.420 66.570 53.345 68.160 ;
        RECT 49.085 64.680 53.345 66.570 ;
        RECT 49.085 64.420 49.515 64.680 ;
        RECT 49.090 64.390 49.510 64.420 ;
        RECT 50.420 63.160 53.345 64.680 ;
        RECT 49.675 62.530 53.345 63.160 ;
        RECT 51.275 61.340 53.345 62.530 ;
        RECT 38.565 30.685 39.515 59.565 ;
        RECT 42.020 54.925 43.215 55.505 ;
        RECT 40.730 54.425 43.215 54.925 ;
        RECT 40.730 54.330 41.150 54.425 ;
        RECT 42.020 54.015 43.215 54.425 ;
        RECT 42.020 51.845 43.215 52.425 ;
        RECT 40.730 51.345 43.215 51.845 ;
        RECT 40.730 51.250 41.150 51.345 ;
        RECT 42.020 50.935 43.215 51.345 ;
        RECT 42.020 48.765 43.215 49.345 ;
        RECT 40.730 48.265 43.215 48.765 ;
        RECT 40.730 48.170 41.150 48.265 ;
        RECT 42.020 47.855 43.215 48.265 ;
        RECT 42.020 45.685 43.215 46.265 ;
        RECT 40.730 45.185 43.215 45.685 ;
        RECT 40.730 45.090 41.150 45.185 ;
        RECT 42.020 44.775 43.215 45.185 ;
        RECT 42.020 42.605 43.215 43.185 ;
        RECT 40.730 42.105 43.215 42.605 ;
        RECT 40.730 42.010 41.150 42.105 ;
        RECT 42.020 41.695 43.215 42.105 ;
        RECT 42.020 39.525 43.215 40.105 ;
        RECT 40.730 39.025 43.215 39.525 ;
        RECT 40.730 38.930 41.150 39.025 ;
        RECT 42.020 38.615 43.215 39.025 ;
        RECT 42.020 36.445 43.215 37.025 ;
        RECT 40.730 35.945 43.215 36.445 ;
        RECT 40.730 35.850 41.150 35.945 ;
        RECT 42.020 35.535 43.215 35.945 ;
        RECT 42.020 33.460 43.215 33.945 ;
        RECT 42.020 33.365 44.545 33.460 ;
        RECT 40.730 32.940 44.545 33.365 ;
        RECT 40.730 32.865 43.215 32.940 ;
        RECT 40.730 32.770 41.150 32.865 ;
        RECT 42.020 32.455 43.215 32.865 ;
        RECT 44.120 32.770 44.540 32.940 ;
        RECT 40.490 21.015 46.255 28.160 ;
        RECT 34.390 20.995 52.780 21.015 ;
        RECT 34.330 20.530 52.840 20.995 ;
        RECT 34.390 20.510 52.780 20.530 ;
        RECT 55.055 20.430 57.215 23.025 ;
      LAYER via ;
        RECT 24.380 80.360 24.640 80.620 ;
        RECT 24.700 80.360 24.960 80.620 ;
        RECT 25.020 80.360 25.280 80.620 ;
        RECT 25.340 80.360 25.600 80.620 ;
        RECT 25.660 80.360 25.920 80.620 ;
        RECT 25.980 80.360 26.240 80.620 ;
        RECT 26.300 80.360 26.560 80.620 ;
        RECT 26.620 80.360 26.880 80.620 ;
        RECT 26.940 80.360 27.200 80.620 ;
        RECT 27.260 80.360 27.520 80.620 ;
        RECT 27.580 80.360 27.840 80.620 ;
        RECT 27.900 80.360 28.160 80.620 ;
        RECT 28.220 80.360 28.480 80.620 ;
        RECT 28.540 80.360 28.800 80.620 ;
        RECT 28.860 80.360 29.120 80.620 ;
        RECT 29.180 80.360 29.440 80.620 ;
        RECT 29.500 80.360 29.760 80.620 ;
        RECT 29.820 80.360 30.080 80.620 ;
        RECT 30.140 80.360 30.400 80.620 ;
        RECT 30.460 80.360 30.720 80.620 ;
        RECT 30.780 80.360 31.040 80.620 ;
        RECT 31.100 80.360 31.360 80.620 ;
        RECT 31.420 80.360 31.680 80.620 ;
        RECT 31.740 80.360 32.000 80.620 ;
        RECT 32.060 80.360 32.320 80.620 ;
        RECT 32.380 80.360 32.640 80.620 ;
        RECT 32.700 80.360 32.960 80.620 ;
        RECT 33.020 80.360 33.280 80.620 ;
        RECT 33.340 80.360 33.600 80.620 ;
        RECT 33.660 80.360 33.920 80.620 ;
        RECT 33.980 80.360 34.240 80.620 ;
        RECT 37.925 76.885 38.185 77.145 ;
        RECT 37.925 76.565 38.185 76.825 ;
        RECT 37.925 76.245 38.185 76.505 ;
        RECT 37.925 75.925 38.185 76.185 ;
        RECT 37.925 75.605 38.185 75.865 ;
        RECT 37.925 75.285 38.185 75.545 ;
        RECT 37.925 74.965 38.185 75.225 ;
        RECT 37.925 74.645 38.185 74.905 ;
        RECT 37.925 74.325 38.185 74.585 ;
        RECT 37.925 74.005 38.185 74.265 ;
        RECT 37.925 73.685 38.185 73.945 ;
        RECT 37.925 73.365 38.185 73.625 ;
        RECT 37.925 73.045 38.185 73.305 ;
        RECT 37.925 72.725 38.185 72.985 ;
        RECT 37.925 72.405 38.185 72.665 ;
        RECT 37.925 72.085 38.185 72.345 ;
        RECT 37.925 71.765 38.185 72.025 ;
        RECT 37.925 71.445 38.185 71.705 ;
        RECT 37.925 71.125 38.185 71.385 ;
        RECT 37.925 70.805 38.185 71.065 ;
        RECT 37.925 70.485 38.185 70.745 ;
        RECT 37.925 70.165 38.185 70.425 ;
        RECT 37.925 69.845 38.185 70.105 ;
        RECT 37.925 69.525 38.185 69.785 ;
        RECT 51.590 61.580 53.130 68.560 ;
        RECT 38.750 59.140 39.010 59.400 ;
        RECT 38.750 58.820 39.010 59.080 ;
        RECT 38.750 58.500 39.010 58.760 ;
        RECT 38.750 58.180 39.010 58.440 ;
        RECT 38.750 57.860 39.010 58.120 ;
        RECT 38.750 57.540 39.010 57.800 ;
        RECT 38.750 57.220 39.010 57.480 ;
        RECT 38.750 56.900 39.010 57.160 ;
        RECT 38.750 56.580 39.010 56.840 ;
        RECT 38.750 56.260 39.010 56.520 ;
        RECT 38.750 55.940 39.010 56.200 ;
        RECT 38.750 55.620 39.010 55.880 ;
        RECT 38.750 55.300 39.010 55.560 ;
        RECT 38.750 54.980 39.010 55.240 ;
        RECT 38.750 54.660 39.010 54.920 ;
        RECT 38.750 54.340 39.010 54.600 ;
        RECT 38.750 54.020 39.010 54.280 ;
        RECT 42.170 54.150 43.070 55.370 ;
        RECT 38.750 53.700 39.010 53.960 ;
        RECT 38.750 53.380 39.010 53.640 ;
        RECT 38.750 53.060 39.010 53.320 ;
        RECT 38.750 52.740 39.010 53.000 ;
        RECT 38.750 52.420 39.010 52.680 ;
        RECT 38.750 52.100 39.010 52.360 ;
        RECT 38.750 51.780 39.010 52.040 ;
        RECT 38.750 51.460 39.010 51.720 ;
        RECT 38.750 51.140 39.010 51.400 ;
        RECT 38.750 50.820 39.010 51.080 ;
        RECT 42.170 51.070 43.070 52.290 ;
        RECT 38.750 50.500 39.010 50.760 ;
        RECT 38.750 50.180 39.010 50.440 ;
        RECT 38.750 49.860 39.010 50.120 ;
        RECT 38.750 49.540 39.010 49.800 ;
        RECT 38.750 49.220 39.010 49.480 ;
        RECT 38.750 48.900 39.010 49.160 ;
        RECT 38.750 48.580 39.010 48.840 ;
        RECT 38.750 48.260 39.010 48.520 ;
        RECT 38.750 47.940 39.010 48.200 ;
        RECT 38.750 47.620 39.010 47.880 ;
        RECT 42.170 47.990 43.070 49.210 ;
        RECT 38.750 47.300 39.010 47.560 ;
        RECT 38.750 46.980 39.010 47.240 ;
        RECT 38.750 46.660 39.010 46.920 ;
        RECT 38.750 46.340 39.010 46.600 ;
        RECT 38.750 46.020 39.010 46.280 ;
        RECT 38.750 45.700 39.010 45.960 ;
        RECT 38.750 45.380 39.010 45.640 ;
        RECT 38.750 45.060 39.010 45.320 ;
        RECT 38.750 44.740 39.010 45.000 ;
        RECT 42.170 44.910 43.070 46.130 ;
        RECT 38.750 44.420 39.010 44.680 ;
        RECT 38.750 44.100 39.010 44.360 ;
        RECT 38.750 43.780 39.010 44.040 ;
        RECT 38.750 43.460 39.010 43.720 ;
        RECT 38.750 43.140 39.010 43.400 ;
        RECT 38.750 42.820 39.010 43.080 ;
        RECT 38.750 42.500 39.010 42.760 ;
        RECT 38.750 42.180 39.010 42.440 ;
        RECT 38.750 41.860 39.010 42.120 ;
        RECT 38.750 41.540 39.010 41.800 ;
        RECT 42.170 41.830 43.070 43.050 ;
        RECT 38.750 41.220 39.010 41.480 ;
        RECT 38.750 40.900 39.010 41.160 ;
        RECT 38.750 40.580 39.010 40.840 ;
        RECT 38.750 40.260 39.010 40.520 ;
        RECT 38.750 39.940 39.010 40.200 ;
        RECT 38.750 39.620 39.010 39.880 ;
        RECT 38.750 39.300 39.010 39.560 ;
        RECT 38.750 38.980 39.010 39.240 ;
        RECT 38.750 38.660 39.010 38.920 ;
        RECT 42.170 38.750 43.070 39.970 ;
        RECT 38.750 38.340 39.010 38.600 ;
        RECT 38.750 38.020 39.010 38.280 ;
        RECT 38.750 37.700 39.010 37.960 ;
        RECT 38.750 37.380 39.010 37.640 ;
        RECT 38.750 37.060 39.010 37.320 ;
        RECT 38.750 36.740 39.010 37.000 ;
        RECT 38.750 36.420 39.010 36.680 ;
        RECT 38.750 36.100 39.010 36.360 ;
        RECT 38.750 35.780 39.010 36.040 ;
        RECT 38.750 35.460 39.010 35.720 ;
        RECT 42.170 35.670 43.070 36.890 ;
        RECT 38.750 35.140 39.010 35.400 ;
        RECT 38.750 34.820 39.010 35.080 ;
        RECT 38.750 34.500 39.010 34.760 ;
        RECT 38.750 34.180 39.010 34.440 ;
        RECT 38.750 33.860 39.010 34.120 ;
        RECT 38.750 33.540 39.010 33.800 ;
        RECT 38.750 33.220 39.010 33.480 ;
        RECT 38.750 32.900 39.010 33.160 ;
        RECT 38.750 32.580 39.010 32.840 ;
        RECT 38.750 32.260 39.010 32.520 ;
        RECT 42.170 32.590 43.070 33.810 ;
        RECT 38.750 31.940 39.010 32.200 ;
        RECT 38.750 31.620 39.010 31.880 ;
        RECT 38.750 31.300 39.010 31.560 ;
        RECT 38.750 30.980 39.010 31.240 ;
        RECT 34.495 20.630 34.755 20.890 ;
        RECT 34.815 20.630 35.075 20.890 ;
        RECT 35.135 20.630 35.395 20.890 ;
        RECT 35.455 20.630 35.715 20.890 ;
        RECT 35.775 20.630 36.035 20.890 ;
        RECT 36.095 20.630 36.355 20.890 ;
        RECT 36.415 20.630 36.675 20.890 ;
        RECT 36.735 20.630 36.995 20.890 ;
        RECT 37.055 20.630 37.315 20.890 ;
        RECT 37.375 20.630 37.635 20.890 ;
        RECT 37.695 20.630 37.955 20.890 ;
        RECT 38.015 20.630 38.275 20.890 ;
        RECT 38.335 20.630 38.595 20.890 ;
        RECT 38.655 20.630 38.915 20.890 ;
        RECT 38.975 20.630 39.235 20.890 ;
        RECT 39.295 20.630 39.555 20.890 ;
        RECT 39.615 20.630 39.875 20.890 ;
        RECT 39.935 20.630 40.195 20.890 ;
        RECT 40.255 20.630 40.515 20.890 ;
        RECT 40.575 20.630 40.835 20.890 ;
        RECT 40.895 20.630 41.155 20.890 ;
        RECT 41.215 20.630 41.475 20.890 ;
        RECT 41.535 20.630 41.795 20.890 ;
        RECT 41.855 20.630 42.115 20.890 ;
        RECT 42.175 20.630 42.435 20.890 ;
        RECT 42.495 20.630 42.755 20.890 ;
        RECT 42.815 20.630 43.075 20.890 ;
        RECT 43.135 20.630 43.395 20.890 ;
        RECT 43.455 20.630 43.715 20.890 ;
        RECT 43.775 20.630 44.035 20.890 ;
        RECT 44.095 20.630 44.355 20.890 ;
        RECT 44.415 20.630 44.675 20.890 ;
        RECT 44.735 20.630 44.995 20.890 ;
        RECT 45.055 20.630 45.315 20.890 ;
        RECT 45.375 20.630 45.635 20.890 ;
        RECT 45.695 20.630 45.955 20.890 ;
        RECT 46.015 20.630 46.275 20.890 ;
        RECT 46.335 20.630 46.595 20.890 ;
        RECT 46.655 20.630 46.915 20.890 ;
        RECT 46.975 20.630 47.235 20.890 ;
        RECT 47.295 20.630 47.555 20.890 ;
        RECT 47.615 20.630 47.875 20.890 ;
        RECT 47.935 20.630 48.195 20.890 ;
        RECT 48.255 20.630 48.515 20.890 ;
        RECT 48.575 20.630 48.835 20.890 ;
        RECT 48.895 20.630 49.155 20.890 ;
        RECT 49.215 20.630 49.475 20.890 ;
        RECT 49.535 20.630 49.795 20.890 ;
        RECT 49.855 20.630 50.115 20.890 ;
        RECT 50.175 20.630 50.435 20.890 ;
        RECT 50.495 20.630 50.755 20.890 ;
        RECT 50.815 20.630 51.075 20.890 ;
        RECT 51.135 20.630 51.395 20.890 ;
        RECT 51.455 20.630 51.715 20.890 ;
        RECT 51.775 20.630 52.035 20.890 ;
        RECT 52.095 20.630 52.355 20.890 ;
        RECT 52.415 20.630 52.675 20.890 ;
        RECT 55.185 20.515 57.045 21.735 ;
      LAYER met2 ;
        RECT 24.330 80.710 34.300 81.210 ;
        RECT 24.325 80.270 34.300 80.710 ;
        RECT 24.330 77.470 34.300 80.270 ;
        RECT 24.330 69.185 38.395 77.470 ;
        RECT 24.330 55.335 34.300 69.185 ;
        RECT 51.275 61.340 53.345 68.750 ;
        RECT 38.480 55.335 39.530 59.770 ;
        RECT 41.810 55.335 43.390 55.830 ;
        RECT 24.330 47.045 43.390 55.335 ;
        RECT 24.330 40.555 34.300 47.045 ;
        RECT 38.480 40.555 39.530 47.045 ;
        RECT 41.810 40.555 43.390 47.045 ;
        RECT 24.330 32.265 43.390 40.555 ;
        RECT 24.330 21.790 34.300 32.265 ;
        RECT 38.480 30.595 39.530 32.265 ;
        RECT 41.810 30.655 43.390 32.265 ;
        RECT 24.330 20.460 57.165 21.790 ;
        RECT 24.330 20.000 34.300 20.460 ;
      LAYER via2 ;
        RECT 27.155 79.735 27.435 80.015 ;
        RECT 27.555 79.735 27.835 80.015 ;
        RECT 27.955 79.735 28.235 80.015 ;
        RECT 28.355 79.735 28.635 80.015 ;
        RECT 30.485 79.735 30.765 80.015 ;
        RECT 30.885 79.735 31.165 80.015 ;
        RECT 31.285 79.735 31.565 80.015 ;
        RECT 31.685 79.735 31.965 80.015 ;
        RECT 27.155 79.140 27.435 79.420 ;
        RECT 27.555 79.140 27.835 79.420 ;
        RECT 27.955 79.140 28.235 79.420 ;
        RECT 28.355 79.140 28.635 79.420 ;
        RECT 30.485 79.140 30.765 79.420 ;
        RECT 30.885 79.140 31.165 79.420 ;
        RECT 31.285 79.140 31.565 79.420 ;
        RECT 31.685 79.140 31.965 79.420 ;
        RECT 27.155 20.635 27.435 20.915 ;
        RECT 27.555 20.635 27.835 20.915 ;
        RECT 27.955 20.635 28.235 20.915 ;
        RECT 28.355 20.635 28.635 20.915 ;
        RECT 30.485 20.635 30.765 20.915 ;
        RECT 30.885 20.635 31.165 20.915 ;
        RECT 31.285 20.635 31.565 20.915 ;
        RECT 31.685 20.635 31.965 20.915 ;
        RECT 27.155 20.040 27.435 20.320 ;
        RECT 27.555 20.040 27.835 20.320 ;
        RECT 27.955 20.040 28.235 20.320 ;
        RECT 28.355 20.040 28.635 20.320 ;
        RECT 30.485 20.040 30.765 20.320 ;
        RECT 30.885 20.040 31.165 20.320 ;
        RECT 31.285 20.040 31.565 20.320 ;
        RECT 31.685 20.040 31.965 20.320 ;
      LAYER met3 ;
        RECT 27.080 79.095 32.080 80.805 ;
        RECT 27.080 19.995 32.080 21.705 ;
      LAYER via3 ;
        RECT 27.135 79.715 27.455 80.035 ;
        RECT 27.535 79.715 27.855 80.035 ;
        RECT 27.935 79.715 28.255 80.035 ;
        RECT 28.335 79.715 28.655 80.035 ;
        RECT 30.465 79.715 30.785 80.035 ;
        RECT 30.865 79.715 31.185 80.035 ;
        RECT 31.265 79.715 31.585 80.035 ;
        RECT 31.665 79.715 31.985 80.035 ;
        RECT 27.135 79.120 27.455 79.440 ;
        RECT 27.535 79.120 27.855 79.440 ;
        RECT 27.935 79.120 28.255 79.440 ;
        RECT 28.335 79.120 28.655 79.440 ;
        RECT 30.465 79.120 30.785 79.440 ;
        RECT 30.865 79.120 31.185 79.440 ;
        RECT 31.265 79.120 31.585 79.440 ;
        RECT 31.665 79.120 31.985 79.440 ;
        RECT 27.135 20.615 27.455 20.935 ;
        RECT 27.535 20.615 27.855 20.935 ;
        RECT 27.935 20.615 28.255 20.935 ;
        RECT 28.335 20.615 28.655 20.935 ;
        RECT 30.465 20.615 30.785 20.935 ;
        RECT 30.865 20.615 31.185 20.935 ;
        RECT 31.265 20.615 31.585 20.935 ;
        RECT 31.665 20.615 31.985 20.935 ;
        RECT 27.135 20.020 27.455 20.340 ;
        RECT 27.535 20.020 27.855 20.340 ;
        RECT 27.935 20.020 28.255 20.340 ;
        RECT 28.335 20.020 28.655 20.340 ;
        RECT 30.465 20.020 30.785 20.340 ;
        RECT 30.865 20.020 31.185 20.340 ;
        RECT 31.265 20.020 31.585 20.340 ;
        RECT 31.665 20.020 31.985 20.340 ;
      LAYER met4 ;
        RECT 27.080 -12.320 32.080 112.960 ;
    END
  END vdda1
  PIN vssa1
    ANTENNADIFFAREA 114.014595 ;
    PORT
      LAYER pwell ;
        RECT 21.025 78.880 37.745 79.310 ;
        RECT 21.025 22.220 21.455 78.880 ;
        RECT 37.315 22.220 37.745 78.880 ;
        RECT 54.275 78.980 70.995 79.410 ;
        RECT 39.545 62.440 40.285 68.470 ;
        RECT 40.995 65.810 43.895 68.490 ;
        RECT 41.005 62.780 43.905 65.460 ;
        RECT 47.215 57.000 50.115 59.680 ;
        RECT 50.215 57.000 53.115 59.680 ;
        RECT 47.205 50.500 50.105 53.180 ;
        RECT 50.205 50.500 53.105 53.180 ;
        RECT 47.205 47.720 50.105 50.400 ;
        RECT 50.205 47.720 53.105 50.400 ;
        RECT 47.205 44.940 50.105 47.620 ;
        RECT 50.205 44.940 53.105 47.620 ;
        RECT 47.205 42.160 50.105 44.840 ;
        RECT 50.205 42.160 53.105 44.840 ;
        RECT 47.205 39.380 50.105 42.060 ;
        RECT 50.205 39.380 53.105 42.060 ;
        RECT 47.205 36.600 50.105 39.280 ;
        RECT 50.205 36.600 53.105 39.280 ;
        RECT 47.205 33.820 50.105 36.500 ;
        RECT 50.205 33.820 53.105 36.500 ;
        RECT 47.205 31.040 50.105 33.720 ;
        RECT 50.205 31.040 53.105 33.720 ;
        RECT 47.215 28.260 50.115 30.940 ;
        RECT 50.205 28.260 53.105 30.940 ;
        RECT 47.215 25.480 50.115 28.160 ;
        RECT 21.025 21.790 37.745 22.220 ;
        RECT 54.275 22.320 54.705 78.980 ;
        RECT 70.565 22.320 70.995 78.980 ;
        RECT 54.275 21.890 70.995 22.320 ;
      LAYER li1 ;
        RECT 20.760 79.010 37.925 79.720 ;
        RECT 20.760 22.090 21.330 79.010 ;
        RECT 37.355 28.180 37.925 79.010 ;
        RECT 53.860 79.110 71.240 79.755 ;
        RECT 38.405 68.300 40.070 68.615 ;
        RECT 38.405 62.610 40.155 68.300 ;
        RECT 40.555 68.110 44.045 68.740 ;
        RECT 40.555 66.170 41.385 68.110 ;
        RECT 42.215 67.460 42.675 67.630 ;
        RECT 43.515 66.170 44.045 68.110 ;
        RECT 40.555 65.090 44.045 66.170 ;
        RECT 40.555 63.160 41.385 65.090 ;
        RECT 42.225 63.640 42.685 63.810 ;
        RECT 43.515 63.160 44.045 65.090 ;
        RECT 38.405 61.595 40.070 62.610 ;
        RECT 40.555 62.530 44.045 63.160 ;
        RECT 46.770 59.525 52.990 60.000 ;
        RECT 46.770 59.385 53.535 59.525 ;
        RECT 46.775 59.320 53.535 59.385 ;
        RECT 46.775 57.360 47.575 59.320 ;
        RECT 49.755 57.360 50.575 59.320 ;
        RECT 51.435 57.860 51.895 58.030 ;
        RECT 52.740 57.360 53.535 59.320 ;
        RECT 46.775 57.190 53.535 57.360 ;
        RECT 46.775 52.990 50.565 57.190 ;
        RECT 52.740 52.990 53.535 57.190 ;
        RECT 46.775 52.820 53.535 52.990 ;
        RECT 46.775 50.860 47.570 52.820 ;
        RECT 49.745 50.860 50.565 52.820 ;
        RECT 51.425 51.360 51.885 51.530 ;
        RECT 52.740 50.860 53.535 52.820 ;
        RECT 46.775 50.690 53.535 50.860 ;
        RECT 46.775 50.210 47.570 50.690 ;
        RECT 49.770 50.210 50.565 50.690 ;
        RECT 52.740 50.210 53.535 50.690 ;
        RECT 46.775 50.040 53.535 50.210 ;
        RECT 46.775 48.080 47.570 50.040 ;
        RECT 49.745 48.080 50.565 50.040 ;
        RECT 51.425 48.580 51.885 48.750 ;
        RECT 52.740 48.080 53.535 50.040 ;
        RECT 46.775 47.910 53.535 48.080 ;
        RECT 46.775 47.430 47.570 47.910 ;
        RECT 49.770 47.430 50.565 47.910 ;
        RECT 52.740 47.430 53.535 47.910 ;
        RECT 46.775 47.260 53.535 47.430 ;
        RECT 46.775 45.300 47.570 47.260 ;
        RECT 49.745 45.300 50.565 47.260 ;
        RECT 51.425 45.800 51.885 45.970 ;
        RECT 52.740 45.300 53.535 47.260 ;
        RECT 46.775 45.130 53.535 45.300 ;
        RECT 46.775 44.650 47.570 45.130 ;
        RECT 49.770 44.650 50.565 45.130 ;
        RECT 52.740 44.650 53.535 45.130 ;
        RECT 46.775 44.480 53.535 44.650 ;
        RECT 46.775 42.520 47.570 44.480 ;
        RECT 49.745 42.520 50.565 44.480 ;
        RECT 51.425 43.020 51.885 43.190 ;
        RECT 52.740 42.520 53.535 44.480 ;
        RECT 46.775 42.350 53.535 42.520 ;
        RECT 46.775 41.870 47.570 42.350 ;
        RECT 49.770 41.870 50.565 42.350 ;
        RECT 52.740 41.870 53.535 42.350 ;
        RECT 46.775 41.700 53.535 41.870 ;
        RECT 46.775 39.740 47.570 41.700 ;
        RECT 49.745 39.740 50.565 41.700 ;
        RECT 51.425 40.240 51.885 40.410 ;
        RECT 52.740 39.740 53.535 41.700 ;
        RECT 46.775 39.570 53.535 39.740 ;
        RECT 46.775 39.090 47.570 39.570 ;
        RECT 49.770 39.090 50.565 39.570 ;
        RECT 52.740 39.090 53.535 39.570 ;
        RECT 46.775 38.920 53.535 39.090 ;
        RECT 46.775 36.960 47.570 38.920 ;
        RECT 49.745 36.960 50.565 38.920 ;
        RECT 51.425 37.460 51.885 37.630 ;
        RECT 52.740 36.960 53.535 38.920 ;
        RECT 46.775 36.790 53.535 36.960 ;
        RECT 46.775 36.310 47.570 36.790 ;
        RECT 49.770 36.310 50.565 36.790 ;
        RECT 52.740 36.310 53.535 36.790 ;
        RECT 46.775 36.140 53.535 36.310 ;
        RECT 46.775 34.180 47.570 36.140 ;
        RECT 49.745 34.180 50.565 36.140 ;
        RECT 51.425 34.680 51.885 34.850 ;
        RECT 52.740 34.180 53.535 36.140 ;
        RECT 46.775 34.010 53.535 34.180 ;
        RECT 46.775 33.530 47.570 34.010 ;
        RECT 49.770 33.530 50.565 34.010 ;
        RECT 52.740 33.530 53.535 34.010 ;
        RECT 46.775 33.360 53.535 33.530 ;
        RECT 46.775 31.400 47.570 33.360 ;
        RECT 49.745 31.400 50.565 33.360 ;
        RECT 51.425 31.900 51.885 32.070 ;
        RECT 52.740 31.400 53.535 33.360 ;
        RECT 46.775 31.230 53.535 31.400 ;
        RECT 46.775 30.750 47.570 31.230 ;
        RECT 49.770 30.750 50.565 31.230 ;
        RECT 52.740 30.750 53.535 31.230 ;
        RECT 46.775 30.580 53.535 30.750 ;
        RECT 46.775 28.620 47.575 30.580 ;
        RECT 49.755 28.620 50.565 30.580 ;
        RECT 51.425 29.120 51.885 29.290 ;
        RECT 52.740 28.620 53.535 30.580 ;
        RECT 46.775 28.450 53.535 28.620 ;
        RECT 37.355 22.480 46.240 28.180 ;
        RECT 46.775 27.970 47.570 28.450 ;
        RECT 49.770 27.970 50.565 28.450 ;
        RECT 46.775 27.800 50.565 27.970 ;
        RECT 46.775 25.840 47.575 27.800 ;
        RECT 48.435 26.340 48.895 26.510 ;
        RECT 49.755 26.390 50.565 27.800 ;
        RECT 49.750 25.840 50.595 26.390 ;
        RECT 46.775 25.610 50.595 25.840 ;
        RECT 52.740 25.655 53.535 28.450 ;
        RECT 46.775 25.100 50.560 25.610 ;
        RECT 37.355 22.090 37.925 22.480 ;
        RECT 20.760 21.475 37.925 22.090 ;
        RECT 53.860 22.190 54.575 79.110 ;
        RECT 70.670 22.190 71.240 79.110 ;
        RECT 53.860 21.530 71.240 22.190 ;
      LAYER mcon ;
        RECT 57.715 79.350 57.885 79.520 ;
        RECT 58.075 79.350 58.245 79.520 ;
        RECT 58.435 79.350 58.605 79.520 ;
        RECT 58.795 79.350 58.965 79.520 ;
        RECT 59.155 79.350 59.325 79.520 ;
        RECT 59.515 79.350 59.685 79.520 ;
        RECT 59.875 79.350 60.045 79.520 ;
        RECT 60.235 79.350 60.405 79.520 ;
        RECT 60.595 79.350 60.765 79.520 ;
        RECT 60.955 79.350 61.125 79.520 ;
        RECT 61.315 79.350 61.485 79.520 ;
        RECT 61.675 79.350 61.845 79.520 ;
        RECT 62.035 79.350 62.205 79.520 ;
        RECT 62.395 79.350 62.565 79.520 ;
        RECT 62.755 79.350 62.925 79.520 ;
        RECT 63.115 79.350 63.285 79.520 ;
        RECT 63.475 79.350 63.645 79.520 ;
        RECT 63.835 79.350 64.005 79.520 ;
        RECT 64.195 79.350 64.365 79.520 ;
        RECT 64.555 79.350 64.725 79.520 ;
        RECT 64.915 79.350 65.085 79.520 ;
        RECT 65.275 79.350 65.445 79.520 ;
        RECT 65.635 79.350 65.805 79.520 ;
        RECT 65.995 79.350 66.165 79.520 ;
        RECT 66.355 79.350 66.525 79.520 ;
        RECT 66.715 79.350 66.885 79.520 ;
        RECT 67.075 79.350 67.245 79.520 ;
        RECT 37.580 68.445 37.750 68.615 ;
        RECT 37.580 68.085 37.750 68.255 ;
        RECT 37.580 67.725 37.750 67.895 ;
        RECT 37.580 67.365 37.750 67.535 ;
        RECT 37.580 67.005 37.750 67.175 ;
        RECT 37.580 66.645 37.750 66.815 ;
        RECT 37.580 66.285 37.750 66.455 ;
        RECT 37.580 65.925 37.750 66.095 ;
        RECT 37.580 65.565 37.750 65.735 ;
        RECT 37.580 65.205 37.750 65.375 ;
        RECT 37.580 64.845 37.750 65.015 ;
        RECT 37.580 64.485 37.750 64.655 ;
        RECT 37.580 64.125 37.750 64.295 ;
        RECT 37.580 63.765 37.750 63.935 ;
        RECT 37.580 63.405 37.750 63.575 ;
        RECT 37.580 63.045 37.750 63.215 ;
        RECT 37.580 62.685 37.750 62.855 ;
        RECT 37.580 62.325 37.750 62.495 ;
        RECT 37.580 61.965 37.750 62.135 ;
        RECT 37.580 61.605 37.750 61.775 ;
        RECT 38.435 61.600 40.045 68.610 ;
        RECT 40.750 67.695 40.920 67.865 ;
        RECT 40.750 67.335 40.920 67.505 ;
        RECT 42.360 67.460 42.530 67.630 ;
        RECT 40.750 66.975 40.920 67.145 ;
        RECT 40.750 66.615 40.920 66.785 ;
        RECT 40.845 65.185 41.735 66.075 ;
        RECT 40.760 64.515 40.930 64.685 ;
        RECT 40.760 64.155 40.930 64.325 ;
        RECT 40.760 63.795 40.930 63.965 ;
        RECT 42.370 63.640 42.540 63.810 ;
        RECT 40.760 63.435 40.930 63.605 ;
        RECT 53.220 59.075 53.390 59.245 ;
        RECT 53.220 58.715 53.390 58.885 ;
        RECT 53.220 58.355 53.390 58.525 ;
        RECT 51.580 57.860 51.750 58.030 ;
        RECT 53.220 57.995 53.390 58.165 ;
        RECT 53.220 57.635 53.390 57.805 ;
        RECT 53.220 57.275 53.390 57.445 ;
        RECT 49.875 54.105 50.405 54.635 ;
        RECT 53.220 56.915 53.390 57.085 ;
        RECT 53.220 56.555 53.390 56.725 ;
        RECT 53.220 56.195 53.390 56.365 ;
        RECT 53.220 55.835 53.390 56.005 ;
        RECT 53.220 55.475 53.390 55.645 ;
        RECT 53.220 55.115 53.390 55.285 ;
        RECT 53.220 54.755 53.390 54.925 ;
        RECT 53.220 54.395 53.390 54.565 ;
        RECT 53.220 54.035 53.390 54.205 ;
        RECT 53.220 53.675 53.390 53.845 ;
        RECT 53.220 53.315 53.390 53.485 ;
        RECT 53.220 52.955 53.390 53.125 ;
        RECT 49.910 50.555 50.440 51.805 ;
        RECT 53.220 52.595 53.390 52.765 ;
        RECT 53.220 52.235 53.390 52.405 ;
        RECT 53.220 51.875 53.390 52.045 ;
        RECT 51.570 51.360 51.740 51.530 ;
        RECT 53.220 51.515 53.390 51.685 ;
        RECT 53.220 51.155 53.390 51.325 ;
        RECT 53.220 50.795 53.390 50.965 ;
        RECT 53.220 50.435 53.390 50.605 ;
        RECT 53.220 50.075 53.390 50.245 ;
        RECT 49.910 47.775 50.440 49.025 ;
        RECT 53.220 49.715 53.390 49.885 ;
        RECT 53.220 49.355 53.390 49.525 ;
        RECT 53.220 48.995 53.390 49.165 ;
        RECT 51.570 48.580 51.740 48.750 ;
        RECT 53.220 48.635 53.390 48.805 ;
        RECT 53.220 48.275 53.390 48.445 ;
        RECT 53.220 47.915 53.390 48.085 ;
        RECT 53.220 47.555 53.390 47.725 ;
        RECT 49.910 44.995 50.440 46.245 ;
        RECT 53.220 47.195 53.390 47.365 ;
        RECT 53.220 46.835 53.390 47.005 ;
        RECT 53.220 46.475 53.390 46.645 ;
        RECT 53.220 46.115 53.390 46.285 ;
        RECT 51.570 45.800 51.740 45.970 ;
        RECT 53.220 45.755 53.390 45.925 ;
        RECT 53.220 45.395 53.390 45.565 ;
        RECT 53.220 45.035 53.390 45.205 ;
        RECT 53.220 44.675 53.390 44.845 ;
        RECT 49.910 42.215 50.440 43.465 ;
        RECT 53.220 44.315 53.390 44.485 ;
        RECT 53.220 43.955 53.390 44.125 ;
        RECT 53.220 43.595 53.390 43.765 ;
        RECT 53.220 43.235 53.390 43.405 ;
        RECT 51.570 43.020 51.740 43.190 ;
        RECT 53.220 42.875 53.390 43.045 ;
        RECT 53.220 42.515 53.390 42.685 ;
        RECT 53.220 42.155 53.390 42.325 ;
        RECT 53.220 41.795 53.390 41.965 ;
        RECT 49.910 39.435 50.440 40.685 ;
        RECT 53.220 41.435 53.390 41.605 ;
        RECT 53.220 41.075 53.390 41.245 ;
        RECT 53.220 40.715 53.390 40.885 ;
        RECT 51.570 40.240 51.740 40.410 ;
        RECT 53.220 40.355 53.390 40.525 ;
        RECT 53.220 39.995 53.390 40.165 ;
        RECT 53.220 39.635 53.390 39.805 ;
        RECT 53.220 39.275 53.390 39.445 ;
        RECT 49.910 36.655 50.440 37.905 ;
        RECT 53.220 38.915 53.390 39.085 ;
        RECT 53.220 38.555 53.390 38.725 ;
        RECT 53.220 38.195 53.390 38.365 ;
        RECT 53.220 37.835 53.390 38.005 ;
        RECT 51.570 37.460 51.740 37.630 ;
        RECT 53.220 37.475 53.390 37.645 ;
        RECT 53.220 37.115 53.390 37.285 ;
        RECT 53.220 36.755 53.390 36.925 ;
        RECT 53.220 36.395 53.390 36.565 ;
        RECT 49.910 33.875 50.440 35.125 ;
        RECT 53.220 36.035 53.390 36.205 ;
        RECT 53.220 35.675 53.390 35.845 ;
        RECT 53.220 35.315 53.390 35.485 ;
        RECT 53.220 34.955 53.390 35.125 ;
        RECT 51.570 34.680 51.740 34.850 ;
        RECT 53.220 34.595 53.390 34.765 ;
        RECT 53.220 34.235 53.390 34.405 ;
        RECT 53.220 33.875 53.390 34.045 ;
        RECT 53.220 33.515 53.390 33.685 ;
        RECT 49.910 31.095 50.440 32.345 ;
        RECT 53.220 33.155 53.390 33.325 ;
        RECT 53.220 32.795 53.390 32.965 ;
        RECT 53.220 32.435 53.390 32.605 ;
        RECT 53.220 32.075 53.390 32.245 ;
        RECT 51.570 31.900 51.740 32.070 ;
        RECT 53.220 31.715 53.390 31.885 ;
        RECT 53.220 31.355 53.390 31.525 ;
        RECT 53.220 30.995 53.390 31.165 ;
        RECT 53.220 30.635 53.390 30.805 ;
        RECT 49.910 28.315 50.440 29.565 ;
        RECT 53.220 30.275 53.390 30.445 ;
        RECT 53.220 29.915 53.390 30.085 ;
        RECT 53.220 29.555 53.390 29.725 ;
        RECT 51.570 29.120 51.740 29.290 ;
        RECT 53.220 29.195 53.390 29.365 ;
        RECT 53.220 28.835 53.390 29.005 ;
        RECT 53.220 28.475 53.390 28.645 ;
        RECT 48.580 26.340 48.750 26.510 ;
        RECT 53.220 28.115 53.390 28.285 ;
        RECT 53.220 27.755 53.390 27.925 ;
        RECT 53.220 27.395 53.390 27.565 ;
        RECT 53.220 27.035 53.390 27.205 ;
        RECT 53.220 26.675 53.390 26.845 ;
        RECT 49.910 25.735 50.440 26.265 ;
        RECT 53.220 26.315 53.390 26.485 ;
        RECT 53.220 25.955 53.390 26.125 ;
        RECT 54.065 54.890 54.235 55.060 ;
        RECT 54.065 54.530 54.235 54.700 ;
        RECT 54.065 54.170 54.235 54.340 ;
        RECT 54.065 53.810 54.235 53.980 ;
        RECT 54.065 53.450 54.235 53.620 ;
        RECT 54.065 53.090 54.235 53.260 ;
        RECT 54.065 52.730 54.235 52.900 ;
        RECT 54.065 52.370 54.235 52.540 ;
        RECT 54.065 52.010 54.235 52.180 ;
        RECT 54.065 51.650 54.235 51.820 ;
        RECT 54.065 51.290 54.235 51.460 ;
        RECT 54.065 50.930 54.235 51.100 ;
        RECT 54.065 50.570 54.235 50.740 ;
        RECT 54.065 50.210 54.235 50.380 ;
        RECT 54.065 49.850 54.235 50.020 ;
        RECT 54.065 49.490 54.235 49.660 ;
        RECT 54.065 49.130 54.235 49.300 ;
        RECT 54.065 48.770 54.235 48.940 ;
        RECT 54.065 48.410 54.235 48.580 ;
        RECT 54.065 48.050 54.235 48.220 ;
        RECT 54.065 47.690 54.235 47.860 ;
        RECT 54.065 47.330 54.235 47.500 ;
        RECT 54.065 46.970 54.235 47.140 ;
        RECT 54.080 37.330 54.250 37.500 ;
        RECT 54.080 36.970 54.250 37.140 ;
        RECT 54.080 36.610 54.250 36.780 ;
        RECT 54.080 36.250 54.250 36.420 ;
        RECT 54.080 35.890 54.250 36.060 ;
        RECT 54.080 35.530 54.250 35.700 ;
        RECT 54.080 35.170 54.250 35.340 ;
        RECT 54.080 34.810 54.250 34.980 ;
        RECT 54.080 34.450 54.250 34.620 ;
        RECT 54.080 34.090 54.250 34.260 ;
        RECT 54.080 33.730 54.250 33.900 ;
        RECT 54.080 33.370 54.250 33.540 ;
        RECT 54.080 33.010 54.250 33.180 ;
        RECT 54.080 32.650 54.250 32.820 ;
        RECT 54.080 32.290 54.250 32.460 ;
        RECT 54.080 31.930 54.250 32.100 ;
        RECT 54.080 31.570 54.250 31.740 ;
        RECT 54.080 31.210 54.250 31.380 ;
        RECT 54.080 30.850 54.250 31.020 ;
        RECT 54.080 30.490 54.250 30.660 ;
        RECT 54.080 30.130 54.250 30.300 ;
        RECT 54.080 29.770 54.250 29.940 ;
        RECT 54.080 29.410 54.250 29.580 ;
        RECT 57.720 21.745 57.890 21.915 ;
        RECT 58.080 21.745 58.250 21.915 ;
        RECT 58.440 21.745 58.610 21.915 ;
        RECT 58.800 21.745 58.970 21.915 ;
        RECT 59.160 21.745 59.330 21.915 ;
        RECT 59.520 21.745 59.690 21.915 ;
        RECT 59.880 21.745 60.050 21.915 ;
        RECT 60.240 21.745 60.410 21.915 ;
        RECT 60.600 21.745 60.770 21.915 ;
        RECT 60.960 21.745 61.130 21.915 ;
        RECT 61.320 21.745 61.490 21.915 ;
        RECT 61.680 21.745 61.850 21.915 ;
        RECT 62.040 21.745 62.210 21.915 ;
        RECT 62.400 21.745 62.570 21.915 ;
        RECT 62.760 21.745 62.930 21.915 ;
        RECT 63.120 21.745 63.290 21.915 ;
        RECT 63.480 21.745 63.650 21.915 ;
        RECT 63.840 21.745 64.010 21.915 ;
        RECT 64.200 21.745 64.370 21.915 ;
        RECT 64.560 21.745 64.730 21.915 ;
        RECT 64.920 21.745 65.090 21.915 ;
        RECT 65.280 21.745 65.450 21.915 ;
        RECT 65.640 21.745 65.810 21.915 ;
        RECT 66.000 21.745 66.170 21.915 ;
        RECT 66.360 21.745 66.530 21.915 ;
        RECT 66.720 21.745 66.890 21.915 ;
        RECT 67.080 21.745 67.250 21.915 ;
      LAYER met1 ;
        RECT 57.575 79.700 67.380 79.720 ;
        RECT 57.515 79.170 67.440 79.700 ;
        RECT 57.575 79.150 67.380 79.170 ;
        RECT 37.355 68.835 38.300 68.840 ;
        RECT 37.355 67.980 40.415 68.835 ;
        RECT 37.355 67.560 42.665 67.980 ;
        RECT 37.355 66.400 41.505 67.560 ;
        RECT 42.235 67.430 42.655 67.560 ;
        RECT 37.355 64.850 41.875 66.400 ;
        RECT 37.355 63.740 41.505 64.850 ;
        RECT 42.245 63.740 42.665 63.840 ;
        RECT 37.355 63.320 42.675 63.740 ;
        RECT 37.355 61.425 40.415 63.320 ;
        RECT 37.405 29.140 38.185 61.425 ;
        RECT 39.415 61.395 40.415 61.425 ;
        RECT 51.455 57.970 51.875 58.060 ;
        RECT 51.440 57.920 51.875 57.970 ;
        RECT 51.435 57.830 51.875 57.920 ;
        RECT 51.435 57.410 51.850 57.830 ;
        RECT 49.655 54.540 50.620 54.790 ;
        RECT 51.435 54.540 51.855 57.410 ;
        RECT 49.655 54.120 51.855 54.540 ;
        RECT 49.655 53.950 50.620 54.120 ;
        RECT 49.740 53.280 50.610 53.950 ;
        RECT 49.750 51.435 50.595 51.880 ;
        RECT 51.445 51.435 51.865 51.560 ;
        RECT 49.750 51.015 51.865 51.435 ;
        RECT 49.750 50.975 50.650 51.015 ;
        RECT 49.750 50.485 50.595 50.975 ;
        RECT 49.750 48.655 50.595 49.100 ;
        RECT 51.445 48.655 51.865 48.780 ;
        RECT 49.750 48.235 51.865 48.655 ;
        RECT 49.750 48.195 50.650 48.235 ;
        RECT 49.750 47.705 50.595 48.195 ;
        RECT 49.750 45.875 50.595 46.320 ;
        RECT 51.445 45.875 51.865 46.000 ;
        RECT 49.750 45.455 51.865 45.875 ;
        RECT 49.750 45.415 50.650 45.455 ;
        RECT 49.750 44.925 50.595 45.415 ;
        RECT 49.750 43.095 50.595 43.540 ;
        RECT 51.445 43.095 51.865 43.220 ;
        RECT 49.750 42.675 51.865 43.095 ;
        RECT 49.750 42.635 50.650 42.675 ;
        RECT 49.750 42.145 50.595 42.635 ;
        RECT 49.750 40.315 50.595 40.760 ;
        RECT 51.445 40.315 51.865 40.440 ;
        RECT 49.750 39.895 51.865 40.315 ;
        RECT 49.750 39.855 50.650 39.895 ;
        RECT 49.750 39.365 50.595 39.855 ;
        RECT 49.750 37.535 50.595 37.980 ;
        RECT 51.445 37.535 51.865 37.660 ;
        RECT 49.750 37.115 51.865 37.535 ;
        RECT 49.750 37.075 50.650 37.115 ;
        RECT 49.750 36.585 50.595 37.075 ;
        RECT 49.750 34.755 50.595 35.200 ;
        RECT 51.445 34.755 51.865 34.880 ;
        RECT 49.750 34.335 51.865 34.755 ;
        RECT 49.750 34.295 50.650 34.335 ;
        RECT 49.750 33.805 50.595 34.295 ;
        RECT 49.750 31.975 50.595 32.420 ;
        RECT 51.445 31.975 51.865 32.100 ;
        RECT 49.750 31.555 51.865 31.975 ;
        RECT 49.750 31.515 50.650 31.555 ;
        RECT 49.750 31.025 50.595 31.515 ;
        RECT 37.390 24.035 38.185 29.140 ;
        RECT 49.750 29.155 50.595 29.640 ;
        RECT 51.445 29.155 51.865 29.320 ;
        RECT 49.750 28.735 51.880 29.155 ;
        RECT 49.750 28.245 50.595 28.735 ;
        RECT 48.455 26.390 48.875 26.540 ;
        RECT 49.750 26.420 50.595 26.440 ;
        RECT 49.690 26.390 50.655 26.420 ;
        RECT 48.450 25.970 50.655 26.390 ;
        RECT 49.690 25.580 50.655 25.970 ;
        RECT 52.740 25.645 53.525 59.515 ;
        RECT 53.920 46.810 54.375 55.225 ;
        RECT 53.935 29.250 54.390 37.665 ;
        RECT 49.750 25.560 50.595 25.580 ;
        RECT 37.390 23.135 38.180 24.035 ;
        RECT 57.580 22.095 67.385 22.115 ;
        RECT 57.520 21.565 67.445 22.095 ;
        RECT 57.580 21.545 67.385 21.565 ;
      LAYER via ;
        RECT 57.710 79.305 57.970 79.565 ;
        RECT 58.030 79.305 58.290 79.565 ;
        RECT 58.350 79.305 58.610 79.565 ;
        RECT 58.670 79.305 58.930 79.565 ;
        RECT 58.990 79.305 59.250 79.565 ;
        RECT 59.310 79.305 59.570 79.565 ;
        RECT 59.630 79.305 59.890 79.565 ;
        RECT 59.950 79.305 60.210 79.565 ;
        RECT 60.270 79.305 60.530 79.565 ;
        RECT 60.590 79.305 60.850 79.565 ;
        RECT 60.910 79.305 61.170 79.565 ;
        RECT 61.230 79.305 61.490 79.565 ;
        RECT 61.550 79.305 61.810 79.565 ;
        RECT 61.870 79.305 62.130 79.565 ;
        RECT 62.190 79.305 62.450 79.565 ;
        RECT 62.510 79.305 62.770 79.565 ;
        RECT 62.830 79.305 63.090 79.565 ;
        RECT 63.150 79.305 63.410 79.565 ;
        RECT 63.470 79.305 63.730 79.565 ;
        RECT 63.790 79.305 64.050 79.565 ;
        RECT 64.110 79.305 64.370 79.565 ;
        RECT 64.430 79.305 64.690 79.565 ;
        RECT 64.750 79.305 65.010 79.565 ;
        RECT 65.070 79.305 65.330 79.565 ;
        RECT 65.390 79.305 65.650 79.565 ;
        RECT 65.710 79.305 65.970 79.565 ;
        RECT 66.030 79.305 66.290 79.565 ;
        RECT 66.350 79.305 66.610 79.565 ;
        RECT 66.670 79.305 66.930 79.565 ;
        RECT 66.990 79.305 67.250 79.565 ;
        RECT 38.470 61.615 40.010 68.595 ;
        RECT 53.175 58.950 53.435 59.210 ;
        RECT 53.175 58.630 53.435 58.890 ;
        RECT 53.175 58.310 53.435 58.570 ;
        RECT 53.175 57.990 53.435 58.250 ;
        RECT 53.175 57.670 53.435 57.930 ;
        RECT 49.885 53.350 50.465 54.570 ;
        RECT 53.175 57.350 53.435 57.610 ;
        RECT 53.175 57.030 53.435 57.290 ;
        RECT 53.175 56.710 53.435 56.970 ;
        RECT 53.175 56.390 53.435 56.650 ;
        RECT 53.175 56.070 53.435 56.330 ;
        RECT 53.175 55.750 53.435 56.010 ;
        RECT 53.175 55.430 53.435 55.690 ;
        RECT 53.175 55.110 53.435 55.370 ;
        RECT 53.175 54.790 53.435 55.050 ;
        RECT 53.175 54.470 53.435 54.730 ;
        RECT 53.175 54.150 53.435 54.410 ;
        RECT 53.175 53.830 53.435 54.090 ;
        RECT 53.175 53.510 53.435 53.770 ;
        RECT 53.175 53.190 53.435 53.450 ;
        RECT 53.175 52.870 53.435 53.130 ;
        RECT 53.175 52.550 53.435 52.810 ;
        RECT 53.175 52.230 53.435 52.490 ;
        RECT 53.175 51.910 53.435 52.170 ;
        RECT 49.885 50.570 50.465 51.790 ;
        RECT 53.175 51.590 53.435 51.850 ;
        RECT 53.175 51.270 53.435 51.530 ;
        RECT 53.175 50.950 53.435 51.210 ;
        RECT 53.175 50.630 53.435 50.890 ;
        RECT 53.175 50.310 53.435 50.570 ;
        RECT 53.175 49.990 53.435 50.250 ;
        RECT 53.175 49.670 53.435 49.930 ;
        RECT 53.175 49.350 53.435 49.610 ;
        RECT 49.885 47.790 50.465 49.010 ;
        RECT 53.175 49.030 53.435 49.290 ;
        RECT 53.175 48.710 53.435 48.970 ;
        RECT 53.175 48.390 53.435 48.650 ;
        RECT 53.175 48.070 53.435 48.330 ;
        RECT 53.175 47.750 53.435 48.010 ;
        RECT 53.175 47.430 53.435 47.690 ;
        RECT 53.175 47.110 53.435 47.370 ;
        RECT 53.175 46.790 53.435 47.050 ;
        RECT 54.020 54.885 54.280 55.145 ;
        RECT 54.020 54.565 54.280 54.825 ;
        RECT 54.020 54.245 54.280 54.505 ;
        RECT 54.020 53.925 54.280 54.185 ;
        RECT 54.020 53.605 54.280 53.865 ;
        RECT 54.020 53.285 54.280 53.545 ;
        RECT 54.020 52.965 54.280 53.225 ;
        RECT 54.020 52.645 54.280 52.905 ;
        RECT 54.020 52.325 54.280 52.585 ;
        RECT 54.020 52.005 54.280 52.265 ;
        RECT 54.020 51.685 54.280 51.945 ;
        RECT 54.020 51.365 54.280 51.625 ;
        RECT 54.020 51.045 54.280 51.305 ;
        RECT 54.020 50.725 54.280 50.985 ;
        RECT 54.020 50.405 54.280 50.665 ;
        RECT 54.020 50.085 54.280 50.345 ;
        RECT 54.020 49.765 54.280 50.025 ;
        RECT 54.020 49.445 54.280 49.705 ;
        RECT 54.020 49.125 54.280 49.385 ;
        RECT 54.020 48.805 54.280 49.065 ;
        RECT 54.020 48.485 54.280 48.745 ;
        RECT 54.020 48.165 54.280 48.425 ;
        RECT 54.020 47.845 54.280 48.105 ;
        RECT 54.020 47.525 54.280 47.785 ;
        RECT 54.020 47.205 54.280 47.465 ;
        RECT 54.020 46.885 54.280 47.145 ;
        RECT 53.175 46.470 53.435 46.730 ;
        RECT 49.885 45.010 50.465 46.230 ;
        RECT 53.175 46.150 53.435 46.410 ;
        RECT 53.175 45.830 53.435 46.090 ;
        RECT 53.175 45.510 53.435 45.770 ;
        RECT 53.175 45.190 53.435 45.450 ;
        RECT 53.175 44.870 53.435 45.130 ;
        RECT 53.175 44.550 53.435 44.810 ;
        RECT 53.175 44.230 53.435 44.490 ;
        RECT 53.175 43.910 53.435 44.170 ;
        RECT 53.175 43.590 53.435 43.850 ;
        RECT 49.885 42.230 50.465 43.450 ;
        RECT 53.175 43.270 53.435 43.530 ;
        RECT 53.175 42.950 53.435 43.210 ;
        RECT 53.175 42.630 53.435 42.890 ;
        RECT 53.175 42.310 53.435 42.570 ;
        RECT 53.175 41.990 53.435 42.250 ;
        RECT 53.175 41.670 53.435 41.930 ;
        RECT 53.175 41.350 53.435 41.610 ;
        RECT 53.175 41.030 53.435 41.290 ;
        RECT 49.885 39.450 50.465 40.670 ;
        RECT 53.175 40.710 53.435 40.970 ;
        RECT 53.175 40.390 53.435 40.650 ;
        RECT 53.175 40.070 53.435 40.330 ;
        RECT 53.175 39.750 53.435 40.010 ;
        RECT 53.175 39.430 53.435 39.690 ;
        RECT 53.175 39.110 53.435 39.370 ;
        RECT 53.175 38.790 53.435 39.050 ;
        RECT 53.175 38.470 53.435 38.730 ;
        RECT 53.175 38.150 53.435 38.410 ;
        RECT 49.885 36.670 50.465 37.890 ;
        RECT 53.175 37.830 53.435 38.090 ;
        RECT 53.175 37.510 53.435 37.770 ;
        RECT 53.175 37.190 53.435 37.450 ;
        RECT 53.175 36.870 53.435 37.130 ;
        RECT 53.175 36.550 53.435 36.810 ;
        RECT 53.175 36.230 53.435 36.490 ;
        RECT 53.175 35.910 53.435 36.170 ;
        RECT 53.175 35.590 53.435 35.850 ;
        RECT 53.175 35.270 53.435 35.530 ;
        RECT 49.885 33.890 50.465 35.110 ;
        RECT 53.175 34.950 53.435 35.210 ;
        RECT 53.175 34.630 53.435 34.890 ;
        RECT 53.175 34.310 53.435 34.570 ;
        RECT 53.175 33.990 53.435 34.250 ;
        RECT 53.175 33.670 53.435 33.930 ;
        RECT 53.175 33.350 53.435 33.610 ;
        RECT 53.175 33.030 53.435 33.290 ;
        RECT 53.175 32.710 53.435 32.970 ;
        RECT 49.885 31.110 50.465 32.330 ;
        RECT 53.175 32.390 53.435 32.650 ;
        RECT 53.175 32.070 53.435 32.330 ;
        RECT 53.175 31.750 53.435 32.010 ;
        RECT 53.175 31.430 53.435 31.690 ;
        RECT 53.175 31.110 53.435 31.370 ;
        RECT 53.175 30.790 53.435 31.050 ;
        RECT 53.175 30.470 53.435 30.730 ;
        RECT 53.175 30.150 53.435 30.410 ;
        RECT 53.175 29.830 53.435 30.090 ;
        RECT 37.490 23.270 38.070 28.970 ;
        RECT 49.885 28.330 50.465 29.550 ;
        RECT 53.175 29.510 53.435 29.770 ;
        RECT 53.175 29.190 53.435 29.450 ;
        RECT 54.035 37.325 54.295 37.585 ;
        RECT 54.035 37.005 54.295 37.265 ;
        RECT 54.035 36.685 54.295 36.945 ;
        RECT 54.035 36.365 54.295 36.625 ;
        RECT 54.035 36.045 54.295 36.305 ;
        RECT 54.035 35.725 54.295 35.985 ;
        RECT 54.035 35.405 54.295 35.665 ;
        RECT 54.035 35.085 54.295 35.345 ;
        RECT 54.035 34.765 54.295 35.025 ;
        RECT 54.035 34.445 54.295 34.705 ;
        RECT 54.035 34.125 54.295 34.385 ;
        RECT 54.035 33.805 54.295 34.065 ;
        RECT 54.035 33.485 54.295 33.745 ;
        RECT 54.035 33.165 54.295 33.425 ;
        RECT 54.035 32.845 54.295 33.105 ;
        RECT 54.035 32.525 54.295 32.785 ;
        RECT 54.035 32.205 54.295 32.465 ;
        RECT 54.035 31.885 54.295 32.145 ;
        RECT 54.035 31.565 54.295 31.825 ;
        RECT 54.035 31.245 54.295 31.505 ;
        RECT 54.035 30.925 54.295 31.185 ;
        RECT 54.035 30.605 54.295 30.865 ;
        RECT 54.035 30.285 54.295 30.545 ;
        RECT 54.035 29.965 54.295 30.225 ;
        RECT 54.035 29.645 54.295 29.905 ;
        RECT 54.035 29.325 54.295 29.585 ;
        RECT 53.175 28.870 53.435 29.130 ;
        RECT 53.175 28.550 53.435 28.810 ;
        RECT 53.175 28.230 53.435 28.490 ;
        RECT 53.175 27.910 53.435 28.170 ;
        RECT 53.175 27.590 53.435 27.850 ;
        RECT 53.175 27.270 53.435 27.530 ;
        RECT 53.175 26.950 53.435 27.210 ;
        RECT 53.175 26.630 53.435 26.890 ;
        RECT 49.885 25.710 50.465 26.290 ;
        RECT 53.175 26.310 53.435 26.570 ;
        RECT 53.175 25.990 53.435 26.250 ;
        RECT 57.715 21.700 57.975 21.960 ;
        RECT 58.035 21.700 58.295 21.960 ;
        RECT 58.355 21.700 58.615 21.960 ;
        RECT 58.675 21.700 58.935 21.960 ;
        RECT 58.995 21.700 59.255 21.960 ;
        RECT 59.315 21.700 59.575 21.960 ;
        RECT 59.635 21.700 59.895 21.960 ;
        RECT 59.955 21.700 60.215 21.960 ;
        RECT 60.275 21.700 60.535 21.960 ;
        RECT 60.595 21.700 60.855 21.960 ;
        RECT 60.915 21.700 61.175 21.960 ;
        RECT 61.235 21.700 61.495 21.960 ;
        RECT 61.555 21.700 61.815 21.960 ;
        RECT 61.875 21.700 62.135 21.960 ;
        RECT 62.195 21.700 62.455 21.960 ;
        RECT 62.515 21.700 62.775 21.960 ;
        RECT 62.835 21.700 63.095 21.960 ;
        RECT 63.155 21.700 63.415 21.960 ;
        RECT 63.475 21.700 63.735 21.960 ;
        RECT 63.795 21.700 64.055 21.960 ;
        RECT 64.115 21.700 64.375 21.960 ;
        RECT 64.435 21.700 64.695 21.960 ;
        RECT 64.755 21.700 65.015 21.960 ;
        RECT 65.075 21.700 65.335 21.960 ;
        RECT 65.395 21.700 65.655 21.960 ;
        RECT 65.715 21.700 65.975 21.960 ;
        RECT 66.035 21.700 66.295 21.960 ;
        RECT 66.355 21.700 66.615 21.960 ;
        RECT 66.675 21.700 66.935 21.960 ;
        RECT 66.995 21.700 67.255 21.960 ;
      LAYER met2 ;
        RECT 37.355 68.835 38.300 68.840 ;
        RECT 37.355 61.425 40.275 68.835 ;
        RECT 49.585 55.170 51.095 55.675 ;
        RECT 52.615 55.170 53.685 59.650 ;
        RECT 57.495 55.170 67.465 81.210 ;
        RECT 49.585 46.875 67.465 55.170 ;
        RECT 49.585 37.600 51.095 46.875 ;
        RECT 52.615 46.870 54.395 46.875 ;
        RECT 52.615 37.605 53.685 46.870 ;
        RECT 52.615 37.600 54.410 37.605 ;
        RECT 57.495 37.600 67.465 46.875 ;
        RECT 49.585 29.305 67.465 37.600 ;
        RECT 37.390 25.875 38.180 29.140 ;
        RECT 40.485 25.875 46.270 28.175 ;
        RECT 49.585 25.875 51.095 29.305 ;
        RECT 52.615 25.875 53.685 29.305 ;
        RECT 57.495 25.875 67.465 29.305 ;
        RECT 37.390 23.135 67.465 25.875 ;
        RECT 37.480 23.125 67.465 23.135 ;
        RECT 57.495 20.000 67.465 23.125 ;
      LAYER via2 ;
        RECT 60.725 79.870 61.005 80.150 ;
        RECT 61.125 79.870 61.405 80.150 ;
        RECT 61.525 79.870 61.805 80.150 ;
        RECT 61.925 79.870 62.205 80.150 ;
        RECT 64.055 79.870 64.335 80.150 ;
        RECT 64.455 79.870 64.735 80.150 ;
        RECT 64.855 79.870 65.135 80.150 ;
        RECT 65.255 79.870 65.535 80.150 ;
        RECT 60.725 79.275 61.005 79.555 ;
        RECT 61.125 79.275 61.405 79.555 ;
        RECT 61.525 79.275 61.805 79.555 ;
        RECT 61.925 79.275 62.205 79.555 ;
        RECT 64.055 79.275 64.335 79.555 ;
        RECT 64.455 79.275 64.735 79.555 ;
        RECT 64.855 79.275 65.135 79.555 ;
        RECT 65.255 79.275 65.535 79.555 ;
        RECT 57.895 35.480 58.975 57.360 ;
        RECT 60.725 20.670 61.005 20.950 ;
        RECT 61.125 20.670 61.405 20.950 ;
        RECT 61.525 20.670 61.805 20.950 ;
        RECT 61.925 20.670 62.205 20.950 ;
        RECT 64.055 20.670 64.335 20.950 ;
        RECT 64.455 20.670 64.735 20.950 ;
        RECT 64.855 20.670 65.135 20.950 ;
        RECT 65.255 20.670 65.535 20.950 ;
        RECT 60.725 20.075 61.005 20.355 ;
        RECT 61.125 20.075 61.405 20.355 ;
        RECT 61.525 20.075 61.805 20.355 ;
        RECT 61.925 20.075 62.205 20.355 ;
        RECT 64.055 20.075 64.335 20.355 ;
        RECT 64.455 20.075 64.735 20.355 ;
        RECT 64.855 20.075 65.135 20.355 ;
        RECT 65.255 20.075 65.535 20.355 ;
      LAYER met3 ;
        RECT 60.650 79.195 65.650 80.905 ;
        RECT 57.740 57.380 59.125 57.435 ;
        RECT 46.750 41.820 53.150 57.340 ;
        RECT 53.700 56.790 59.125 57.380 ;
        RECT 57.740 52.050 59.125 56.790 ;
        RECT 53.700 51.460 59.125 52.050 ;
        RECT 57.740 46.720 59.125 51.460 ;
        RECT 53.700 46.130 59.125 46.720 ;
        RECT 46.755 31.160 53.155 41.820 ;
        RECT 57.740 41.390 59.125 46.130 ;
        RECT 53.700 40.800 59.125 41.390 ;
        RECT 57.740 36.060 59.125 40.800 ;
        RECT 53.700 35.470 59.125 36.060 ;
        RECT 57.740 35.405 59.125 35.470 ;
        RECT 60.650 19.995 65.650 21.705 ;
      LAYER via3 ;
        RECT 60.705 79.850 61.025 80.170 ;
        RECT 61.105 79.850 61.425 80.170 ;
        RECT 61.505 79.850 61.825 80.170 ;
        RECT 61.905 79.850 62.225 80.170 ;
        RECT 64.035 79.850 64.355 80.170 ;
        RECT 64.435 79.850 64.755 80.170 ;
        RECT 64.835 79.850 65.155 80.170 ;
        RECT 65.235 79.850 65.555 80.170 ;
        RECT 60.705 79.255 61.025 79.575 ;
        RECT 61.105 79.255 61.425 79.575 ;
        RECT 61.505 79.255 61.825 79.575 ;
        RECT 61.905 79.255 62.225 79.575 ;
        RECT 64.035 79.255 64.355 79.575 ;
        RECT 64.435 79.255 64.755 79.575 ;
        RECT 64.835 79.255 65.155 79.575 ;
        RECT 65.235 79.255 65.555 79.575 ;
        RECT 46.990 56.920 47.310 57.240 ;
        RECT 47.390 56.920 47.710 57.240 ;
        RECT 47.790 56.920 48.110 57.240 ;
        RECT 48.190 56.920 48.510 57.240 ;
        RECT 48.590 56.920 48.910 57.240 ;
        RECT 48.990 56.920 49.310 57.240 ;
        RECT 49.390 56.920 49.710 57.240 ;
        RECT 49.790 56.920 50.110 57.240 ;
        RECT 50.190 56.920 50.510 57.240 ;
        RECT 50.590 56.920 50.910 57.240 ;
        RECT 50.990 56.920 51.310 57.240 ;
        RECT 51.390 56.920 51.710 57.240 ;
        RECT 51.790 56.920 52.110 57.240 ;
        RECT 52.190 56.920 52.510 57.240 ;
        RECT 52.590 56.920 52.910 57.240 ;
        RECT 53.765 56.925 54.085 57.245 ;
        RECT 54.165 56.925 54.485 57.245 ;
        RECT 54.565 56.925 54.885 57.245 ;
        RECT 46.990 51.590 47.310 51.910 ;
        RECT 47.390 51.590 47.710 51.910 ;
        RECT 47.790 51.590 48.110 51.910 ;
        RECT 48.190 51.590 48.510 51.910 ;
        RECT 48.590 51.590 48.910 51.910 ;
        RECT 48.990 51.590 49.310 51.910 ;
        RECT 49.390 51.590 49.710 51.910 ;
        RECT 49.790 51.590 50.110 51.910 ;
        RECT 50.190 51.590 50.510 51.910 ;
        RECT 50.590 51.590 50.910 51.910 ;
        RECT 50.990 51.590 51.310 51.910 ;
        RECT 51.390 51.590 51.710 51.910 ;
        RECT 51.790 51.590 52.110 51.910 ;
        RECT 52.190 51.590 52.510 51.910 ;
        RECT 52.590 51.590 52.910 51.910 ;
        RECT 53.765 51.595 54.085 51.915 ;
        RECT 54.165 51.595 54.485 51.915 ;
        RECT 54.565 51.595 54.885 51.915 ;
        RECT 46.990 46.260 47.310 46.580 ;
        RECT 47.390 46.260 47.710 46.580 ;
        RECT 47.790 46.260 48.110 46.580 ;
        RECT 48.190 46.260 48.510 46.580 ;
        RECT 48.590 46.260 48.910 46.580 ;
        RECT 48.990 46.260 49.310 46.580 ;
        RECT 49.390 46.260 49.710 46.580 ;
        RECT 49.790 46.260 50.110 46.580 ;
        RECT 50.190 46.260 50.510 46.580 ;
        RECT 50.590 46.260 50.910 46.580 ;
        RECT 50.990 46.260 51.310 46.580 ;
        RECT 51.390 46.260 51.710 46.580 ;
        RECT 51.790 46.260 52.110 46.580 ;
        RECT 52.190 46.260 52.510 46.580 ;
        RECT 52.590 46.260 52.910 46.580 ;
        RECT 53.765 46.265 54.085 46.585 ;
        RECT 54.165 46.265 54.485 46.585 ;
        RECT 54.565 46.265 54.885 46.585 ;
        RECT 46.995 40.930 47.315 41.250 ;
        RECT 47.395 40.930 47.715 41.250 ;
        RECT 47.795 40.930 48.115 41.250 ;
        RECT 48.195 40.930 48.515 41.250 ;
        RECT 48.595 40.930 48.915 41.250 ;
        RECT 48.995 40.930 49.315 41.250 ;
        RECT 49.395 40.930 49.715 41.250 ;
        RECT 49.795 40.930 50.115 41.250 ;
        RECT 50.195 40.930 50.515 41.250 ;
        RECT 50.595 40.930 50.915 41.250 ;
        RECT 50.995 40.930 51.315 41.250 ;
        RECT 51.395 40.930 51.715 41.250 ;
        RECT 51.795 40.930 52.115 41.250 ;
        RECT 52.195 40.930 52.515 41.250 ;
        RECT 52.595 40.930 52.915 41.250 ;
        RECT 53.765 40.935 54.085 41.255 ;
        RECT 54.165 40.935 54.485 41.255 ;
        RECT 54.565 40.935 54.885 41.255 ;
        RECT 46.995 35.600 47.315 35.920 ;
        RECT 47.395 35.600 47.715 35.920 ;
        RECT 47.795 35.600 48.115 35.920 ;
        RECT 48.195 35.600 48.515 35.920 ;
        RECT 48.595 35.600 48.915 35.920 ;
        RECT 48.995 35.600 49.315 35.920 ;
        RECT 49.395 35.600 49.715 35.920 ;
        RECT 49.795 35.600 50.115 35.920 ;
        RECT 50.195 35.600 50.515 35.920 ;
        RECT 50.595 35.600 50.915 35.920 ;
        RECT 50.995 35.600 51.315 35.920 ;
        RECT 51.395 35.600 51.715 35.920 ;
        RECT 51.795 35.600 52.115 35.920 ;
        RECT 52.195 35.600 52.515 35.920 ;
        RECT 52.595 35.600 52.915 35.920 ;
        RECT 53.765 35.605 54.085 35.925 ;
        RECT 54.165 35.605 54.485 35.925 ;
        RECT 54.565 35.605 54.885 35.925 ;
        RECT 60.705 20.650 61.025 20.970 ;
        RECT 61.105 20.650 61.425 20.970 ;
        RECT 61.505 20.650 61.825 20.970 ;
        RECT 61.905 20.650 62.225 20.970 ;
        RECT 64.035 20.650 64.355 20.970 ;
        RECT 64.435 20.650 64.755 20.970 ;
        RECT 64.835 20.650 65.155 20.970 ;
        RECT 65.235 20.650 65.555 20.970 ;
        RECT 60.705 20.055 61.025 20.375 ;
        RECT 61.105 20.055 61.425 20.375 ;
        RECT 61.505 20.055 61.825 20.375 ;
        RECT 61.905 20.055 62.225 20.375 ;
        RECT 64.035 20.055 64.355 20.375 ;
        RECT 64.435 20.055 64.755 20.375 ;
        RECT 64.835 20.055 65.155 20.375 ;
        RECT 65.235 20.055 65.555 20.375 ;
      LAYER met4 ;
        RECT 53.695 57.330 54.955 57.335 ;
        RECT 52.405 57.320 54.955 57.330 ;
        RECT 46.810 56.840 54.955 57.320 ;
        RECT 53.695 56.835 54.955 56.840 ;
        RECT 53.695 52.000 54.955 52.005 ;
        RECT 52.405 51.990 54.955 52.000 ;
        RECT 46.810 51.510 54.955 51.990 ;
        RECT 53.695 51.505 54.955 51.510 ;
        RECT 53.695 46.670 54.955 46.675 ;
        RECT 52.405 46.660 54.955 46.670 ;
        RECT 46.810 46.180 54.955 46.660 ;
        RECT 53.695 46.175 54.955 46.180 ;
        RECT 53.695 41.340 54.955 41.345 ;
        RECT 52.405 41.330 54.955 41.340 ;
        RECT 46.815 40.850 54.955 41.330 ;
        RECT 53.695 40.845 54.955 40.850 ;
        RECT 53.695 36.010 54.955 36.015 ;
        RECT 52.405 36.000 54.955 36.010 ;
        RECT 46.815 35.520 54.955 36.000 ;
        RECT 53.695 35.515 54.955 35.520 ;
        RECT 60.650 -12.320 65.650 112.960 ;
    END
  END vssa1
  OBS
      LAYER li1 ;
        RECT 42.590 79.510 43.130 79.680 ;
        RECT 43.300 79.210 43.470 79.540 ;
        RECT 45.455 79.225 45.625 79.555 ;
        RECT 48.410 79.545 48.950 79.715 ;
        RECT 21.805 78.180 23.965 78.530 ;
        RECT 34.805 78.180 36.965 78.530 ;
        RECT 55.055 78.280 57.215 78.630 ;
        RECT 68.055 78.280 70.215 78.630 ;
        RECT 21.805 77.350 23.965 77.700 ;
        RECT 34.805 77.350 36.965 77.700 ;
        RECT 55.055 77.450 57.215 77.800 ;
        RECT 68.055 77.450 70.215 77.800 ;
        RECT 21.805 76.520 23.965 76.870 ;
        RECT 34.805 76.520 36.965 76.870 ;
        RECT 46.670 76.705 47.130 76.875 ;
        RECT 55.055 76.620 57.215 76.970 ;
        RECT 68.055 76.620 70.215 76.970 ;
        RECT 21.805 75.690 23.965 76.040 ;
        RECT 34.805 75.690 36.965 76.040 ;
        RECT 55.055 75.790 57.215 76.140 ;
        RECT 68.055 75.790 70.215 76.140 ;
        RECT 21.805 74.860 23.965 75.210 ;
        RECT 34.805 74.860 36.965 75.210 ;
        RECT 43.545 75.120 44.585 75.290 ;
        RECT 46.735 75.120 47.775 75.290 ;
        RECT 55.055 74.960 57.215 75.310 ;
        RECT 68.055 74.960 70.215 75.310 ;
        RECT 21.805 74.030 23.965 74.380 ;
        RECT 34.805 74.030 36.965 74.380 ;
        RECT 55.055 74.130 57.215 74.480 ;
        RECT 68.055 74.130 70.215 74.480 ;
        RECT 21.805 73.200 23.965 73.550 ;
        RECT 34.805 73.200 36.965 73.550 ;
        RECT 55.055 73.300 57.215 73.650 ;
        RECT 68.055 73.300 70.215 73.650 ;
        RECT 21.805 72.370 23.965 72.720 ;
        RECT 34.805 72.370 36.965 72.720 ;
        RECT 55.055 72.470 57.215 72.820 ;
        RECT 68.055 72.470 70.215 72.820 ;
        RECT 21.805 71.540 23.965 71.890 ;
        RECT 34.805 71.540 36.965 71.890 ;
        RECT 42.485 71.670 42.655 72.000 ;
        RECT 55.055 71.640 57.215 71.990 ;
        RECT 68.055 71.640 70.215 71.990 ;
        RECT 21.805 70.710 23.965 71.060 ;
        RECT 34.805 70.710 36.965 71.060 ;
        RECT 55.055 70.810 57.215 71.160 ;
        RECT 68.055 70.810 70.215 71.160 ;
        RECT 21.805 69.880 23.965 70.230 ;
        RECT 34.805 69.880 36.965 70.230 ;
        RECT 55.055 69.980 57.215 70.330 ;
        RECT 68.055 69.980 70.215 70.330 ;
        RECT 21.805 69.050 23.965 69.400 ;
        RECT 34.805 69.050 36.965 69.400 ;
        RECT 55.055 69.150 57.215 69.500 ;
        RECT 68.055 69.150 70.215 69.500 ;
        RECT 21.805 68.220 23.965 68.570 ;
        RECT 34.805 68.220 36.965 68.570 ;
        RECT 55.055 68.320 57.215 68.670 ;
        RECT 68.055 68.320 70.215 68.670 ;
        RECT 21.805 67.390 23.965 67.740 ;
        RECT 34.805 67.390 36.965 67.740 ;
        RECT 45.730 67.470 46.190 67.640 ;
        RECT 49.070 67.500 49.530 67.670 ;
        RECT 55.055 67.490 57.215 67.840 ;
        RECT 68.055 67.490 70.215 67.840 ;
        RECT 45.345 66.910 45.515 67.410 ;
        RECT 46.405 66.910 46.575 67.410 ;
        RECT 48.685 66.940 48.855 67.440 ;
        RECT 49.745 66.940 49.915 67.440 ;
        RECT 21.805 66.560 23.965 66.910 ;
        RECT 34.805 66.560 36.965 66.910 ;
        RECT 42.215 66.670 42.675 66.840 ;
        RECT 45.730 66.680 46.190 66.850 ;
        RECT 55.055 66.660 57.215 67.010 ;
        RECT 68.055 66.660 70.215 67.010 ;
        RECT 21.805 65.730 23.965 66.080 ;
        RECT 34.805 65.730 36.965 66.080 ;
        RECT 55.055 65.830 57.215 66.180 ;
        RECT 68.055 65.830 70.215 66.180 ;
        RECT 21.805 64.900 23.965 65.250 ;
        RECT 34.805 64.900 36.965 65.250 ;
        RECT 55.055 65.000 57.215 65.350 ;
        RECT 68.055 65.000 70.215 65.350 ;
        RECT 42.225 64.430 42.685 64.600 ;
        RECT 45.720 64.420 46.180 64.590 ;
        RECT 21.805 64.070 23.965 64.420 ;
        RECT 34.805 64.070 36.965 64.420 ;
        RECT 41.885 63.870 42.055 64.370 ;
        RECT 42.855 63.870 43.025 64.370 ;
        RECT 45.335 63.860 45.505 64.360 ;
        RECT 46.395 63.860 46.565 64.360 ;
        RECT 48.685 63.860 48.855 64.360 ;
        RECT 49.745 63.860 49.915 64.360 ;
        RECT 55.055 64.170 57.215 64.520 ;
        RECT 68.055 64.170 70.215 64.520 ;
        RECT 45.720 63.630 46.180 63.800 ;
        RECT 49.070 63.630 49.530 63.800 ;
        RECT 21.805 63.240 23.965 63.590 ;
        RECT 34.805 63.240 36.965 63.590 ;
        RECT 55.055 63.340 57.215 63.690 ;
        RECT 68.055 63.340 70.215 63.690 ;
        RECT 21.805 62.410 23.965 62.760 ;
        RECT 34.805 62.410 36.965 62.760 ;
        RECT 55.055 62.510 57.215 62.860 ;
        RECT 68.055 62.510 70.215 62.860 ;
        RECT 21.805 61.580 23.965 61.930 ;
        RECT 34.805 61.580 36.965 61.930 ;
        RECT 55.055 61.680 57.215 62.030 ;
        RECT 68.055 61.680 70.215 62.030 ;
        RECT 21.805 60.750 23.965 61.100 ;
        RECT 34.805 60.750 36.965 61.100 ;
        RECT 55.055 60.850 57.215 61.200 ;
        RECT 68.055 60.850 70.215 61.200 ;
        RECT 21.805 59.920 23.965 60.270 ;
        RECT 34.805 59.920 36.965 60.270 ;
        RECT 55.055 60.020 57.215 60.370 ;
        RECT 68.055 60.020 70.215 60.370 ;
        RECT 21.805 59.090 23.965 59.440 ;
        RECT 34.805 59.090 36.965 59.440 ;
        RECT 55.055 59.190 57.215 59.540 ;
        RECT 68.055 59.190 70.215 59.540 ;
        RECT 44.100 58.710 44.560 58.880 ;
        RECT 48.435 58.650 48.895 58.820 ;
        RECT 51.435 58.650 51.895 58.820 ;
        RECT 21.805 58.260 23.965 58.610 ;
        RECT 34.805 58.260 36.965 58.610 ;
        RECT 43.715 58.150 43.885 58.650 ;
        RECT 44.775 58.150 44.945 58.650 ;
        RECT 51.095 58.090 51.265 58.590 ;
        RECT 52.065 58.090 52.235 58.590 ;
        RECT 55.055 58.360 57.215 58.710 ;
        RECT 68.055 58.360 70.215 58.710 ;
        RECT 48.435 57.860 48.895 58.030 ;
        RECT 21.805 57.430 23.965 57.780 ;
        RECT 34.805 57.430 36.965 57.780 ;
        RECT 55.055 57.530 57.215 57.880 ;
        RECT 68.055 57.530 70.215 57.880 ;
        RECT 21.805 56.600 23.965 56.950 ;
        RECT 34.805 56.600 36.965 56.950 ;
        RECT 55.055 56.700 57.215 57.050 ;
        RECT 68.055 56.700 70.215 57.050 ;
        RECT 21.805 55.770 23.965 56.120 ;
        RECT 34.805 55.770 36.965 56.120 ;
        RECT 55.055 55.870 57.215 56.220 ;
        RECT 68.055 55.870 70.215 56.220 ;
        RECT 21.805 54.940 23.965 55.290 ;
        RECT 34.805 54.940 36.965 55.290 ;
        RECT 55.055 55.040 57.215 55.390 ;
        RECT 68.055 55.040 70.215 55.390 ;
        RECT 21.805 54.110 23.965 54.460 ;
        RECT 34.805 54.110 36.965 54.460 ;
        RECT 44.100 54.360 44.560 54.530 ;
        RECT 40.325 53.800 40.495 54.300 ;
        RECT 41.385 53.800 41.555 54.300 ;
        RECT 43.715 53.800 43.885 54.300 ;
        RECT 44.775 53.800 44.945 54.300 ;
        RECT 55.055 54.210 57.215 54.560 ;
        RECT 68.055 54.210 70.215 54.560 ;
        RECT 21.805 53.280 23.965 53.630 ;
        RECT 34.805 53.280 36.965 53.630 ;
        RECT 40.710 53.570 41.170 53.740 ;
        RECT 44.100 53.570 44.560 53.740 ;
        RECT 55.055 53.380 57.215 53.730 ;
        RECT 68.055 53.380 70.215 53.730 ;
        RECT 21.805 52.450 23.965 52.800 ;
        RECT 34.805 52.450 36.965 52.800 ;
        RECT 55.055 52.550 57.215 52.900 ;
        RECT 68.055 52.550 70.215 52.900 ;
        RECT 48.425 52.150 48.885 52.320 ;
        RECT 51.425 52.150 51.885 52.320 ;
        RECT 21.805 51.620 23.965 51.970 ;
        RECT 34.805 51.620 36.965 51.970 ;
        RECT 48.085 51.590 48.255 52.090 ;
        RECT 49.055 51.590 49.225 52.090 ;
        RECT 51.085 51.590 51.255 52.090 ;
        RECT 52.055 51.590 52.225 52.090 ;
        RECT 55.055 51.720 57.215 52.070 ;
        RECT 68.055 51.720 70.215 52.070 ;
        RECT 44.100 51.280 44.560 51.450 ;
        RECT 48.425 51.360 48.885 51.530 ;
        RECT 21.805 50.790 23.965 51.140 ;
        RECT 34.805 50.790 36.965 51.140 ;
        RECT 40.325 50.720 40.495 51.220 ;
        RECT 41.385 50.720 41.555 51.220 ;
        RECT 43.715 50.720 43.885 51.220 ;
        RECT 44.775 50.720 44.945 51.220 ;
        RECT 55.055 50.890 57.215 51.240 ;
        RECT 68.055 50.890 70.215 51.240 ;
        RECT 40.710 50.490 41.170 50.660 ;
        RECT 44.100 50.490 44.560 50.660 ;
        RECT 21.805 49.960 23.965 50.310 ;
        RECT 34.805 49.960 36.965 50.310 ;
        RECT 55.055 50.060 57.215 50.410 ;
        RECT 68.055 50.060 70.215 50.410 ;
        RECT 21.805 49.130 23.965 49.480 ;
        RECT 34.805 49.130 36.965 49.480 ;
        RECT 48.425 49.370 48.885 49.540 ;
        RECT 51.425 49.370 51.885 49.540 ;
        RECT 48.085 48.810 48.255 49.310 ;
        RECT 49.055 48.810 49.225 49.310 ;
        RECT 51.085 48.810 51.255 49.310 ;
        RECT 52.055 48.810 52.225 49.310 ;
        RECT 55.055 49.230 57.215 49.580 ;
        RECT 68.055 49.230 70.215 49.580 ;
        RECT 21.805 48.300 23.965 48.650 ;
        RECT 34.805 48.300 36.965 48.650 ;
        RECT 48.425 48.580 48.885 48.750 ;
        RECT 55.055 48.400 57.215 48.750 ;
        RECT 68.055 48.400 70.215 48.750 ;
        RECT 44.100 48.200 44.560 48.370 ;
        RECT 21.805 47.470 23.965 47.820 ;
        RECT 34.805 47.470 36.965 47.820 ;
        RECT 40.325 47.640 40.495 48.140 ;
        RECT 41.385 47.640 41.555 48.140 ;
        RECT 43.715 47.640 43.885 48.140 ;
        RECT 44.775 47.640 44.945 48.140 ;
        RECT 40.710 47.410 41.170 47.580 ;
        RECT 44.100 47.410 44.560 47.580 ;
        RECT 55.055 47.570 57.215 47.920 ;
        RECT 68.055 47.570 70.215 47.920 ;
        RECT 21.805 46.640 23.965 46.990 ;
        RECT 34.805 46.640 36.965 46.990 ;
        RECT 48.425 46.590 48.885 46.760 ;
        RECT 51.425 46.590 51.885 46.760 ;
        RECT 55.055 46.740 57.215 47.090 ;
        RECT 68.055 46.740 70.215 47.090 ;
        RECT 21.805 45.810 23.965 46.160 ;
        RECT 34.805 45.810 36.965 46.160 ;
        RECT 48.085 46.030 48.255 46.530 ;
        RECT 49.055 46.030 49.225 46.530 ;
        RECT 51.085 46.030 51.255 46.530 ;
        RECT 52.055 46.030 52.225 46.530 ;
        RECT 48.425 45.800 48.885 45.970 ;
        RECT 55.055 45.910 57.215 46.260 ;
        RECT 68.055 45.910 70.215 46.260 ;
        RECT 21.805 44.980 23.965 45.330 ;
        RECT 34.805 44.980 36.965 45.330 ;
        RECT 44.100 45.120 44.560 45.290 ;
        RECT 55.055 45.080 57.215 45.430 ;
        RECT 68.055 45.080 70.215 45.430 ;
        RECT 40.325 44.560 40.495 45.060 ;
        RECT 41.385 44.560 41.555 45.060 ;
        RECT 43.715 44.560 43.885 45.060 ;
        RECT 44.775 44.560 44.945 45.060 ;
        RECT 21.805 44.150 23.965 44.500 ;
        RECT 34.805 44.150 36.965 44.500 ;
        RECT 40.710 44.330 41.170 44.500 ;
        RECT 44.100 44.330 44.560 44.500 ;
        RECT 55.055 44.250 57.215 44.600 ;
        RECT 68.055 44.250 70.215 44.600 ;
        RECT 48.425 43.810 48.885 43.980 ;
        RECT 51.425 43.810 51.885 43.980 ;
        RECT 21.805 43.320 23.965 43.670 ;
        RECT 34.805 43.320 36.965 43.670 ;
        RECT 48.085 43.250 48.255 43.750 ;
        RECT 49.055 43.250 49.225 43.750 ;
        RECT 51.085 43.250 51.255 43.750 ;
        RECT 52.055 43.250 52.225 43.750 ;
        RECT 55.055 43.420 57.215 43.770 ;
        RECT 68.055 43.420 70.215 43.770 ;
        RECT 48.425 43.020 48.885 43.190 ;
        RECT 21.805 42.490 23.965 42.840 ;
        RECT 34.805 42.490 36.965 42.840 ;
        RECT 55.055 42.590 57.215 42.940 ;
        RECT 68.055 42.590 70.215 42.940 ;
        RECT 44.100 42.040 44.560 42.210 ;
        RECT 21.805 41.660 23.965 42.010 ;
        RECT 34.805 41.660 36.965 42.010 ;
        RECT 40.325 41.480 40.495 41.980 ;
        RECT 41.385 41.480 41.555 41.980 ;
        RECT 43.715 41.480 43.885 41.980 ;
        RECT 44.775 41.480 44.945 41.980 ;
        RECT 55.055 41.760 57.215 42.110 ;
        RECT 68.055 41.760 70.215 42.110 ;
        RECT 40.710 41.250 41.170 41.420 ;
        RECT 44.100 41.250 44.560 41.420 ;
        RECT 21.805 40.830 23.965 41.180 ;
        RECT 34.805 40.830 36.965 41.180 ;
        RECT 48.425 41.030 48.885 41.200 ;
        RECT 51.425 41.030 51.885 41.200 ;
        RECT 48.085 40.470 48.255 40.970 ;
        RECT 49.055 40.470 49.225 40.970 ;
        RECT 51.085 40.470 51.255 40.970 ;
        RECT 52.055 40.470 52.225 40.970 ;
        RECT 55.055 40.930 57.215 41.280 ;
        RECT 68.055 40.930 70.215 41.280 ;
        RECT 21.805 40.000 23.965 40.350 ;
        RECT 34.805 40.000 36.965 40.350 ;
        RECT 48.425 40.240 48.885 40.410 ;
        RECT 55.055 40.100 57.215 40.450 ;
        RECT 68.055 40.100 70.215 40.450 ;
        RECT 21.805 39.170 23.965 39.520 ;
        RECT 34.805 39.170 36.965 39.520 ;
        RECT 55.055 39.270 57.215 39.620 ;
        RECT 68.055 39.270 70.215 39.620 ;
        RECT 44.100 38.960 44.560 39.130 ;
        RECT 21.805 38.340 23.965 38.690 ;
        RECT 34.805 38.340 36.965 38.690 ;
        RECT 40.325 38.400 40.495 38.900 ;
        RECT 41.385 38.400 41.555 38.900 ;
        RECT 43.715 38.400 43.885 38.900 ;
        RECT 44.775 38.400 44.945 38.900 ;
        RECT 55.055 38.440 57.215 38.790 ;
        RECT 68.055 38.440 70.215 38.790 ;
        RECT 40.710 38.170 41.170 38.340 ;
        RECT 44.100 38.170 44.560 38.340 ;
        RECT 48.425 38.250 48.885 38.420 ;
        RECT 51.425 38.250 51.885 38.420 ;
        RECT 21.805 37.510 23.965 37.860 ;
        RECT 34.805 37.510 36.965 37.860 ;
        RECT 48.085 37.690 48.255 38.190 ;
        RECT 49.055 37.690 49.225 38.190 ;
        RECT 51.085 37.690 51.255 38.190 ;
        RECT 52.055 37.690 52.225 38.190 ;
        RECT 48.425 37.460 48.885 37.630 ;
        RECT 55.055 37.610 57.215 37.960 ;
        RECT 68.055 37.610 70.215 37.960 ;
        RECT 21.805 36.680 23.965 37.030 ;
        RECT 34.805 36.680 36.965 37.030 ;
        RECT 55.055 36.780 57.215 37.130 ;
        RECT 68.055 36.780 70.215 37.130 ;
        RECT 21.805 35.850 23.965 36.200 ;
        RECT 34.805 35.850 36.965 36.200 ;
        RECT 44.100 35.880 44.560 36.050 ;
        RECT 55.055 35.950 57.215 36.300 ;
        RECT 68.055 35.950 70.215 36.300 ;
        RECT 21.805 35.020 23.965 35.370 ;
        RECT 34.805 35.020 36.965 35.370 ;
        RECT 40.325 35.320 40.495 35.820 ;
        RECT 41.385 35.320 41.555 35.820 ;
        RECT 43.715 35.320 43.885 35.820 ;
        RECT 44.775 35.320 44.945 35.820 ;
        RECT 48.425 35.470 48.885 35.640 ;
        RECT 51.425 35.470 51.885 35.640 ;
        RECT 40.710 35.090 41.170 35.260 ;
        RECT 44.100 35.090 44.560 35.260 ;
        RECT 48.085 34.910 48.255 35.410 ;
        RECT 49.055 34.910 49.225 35.410 ;
        RECT 51.085 34.910 51.255 35.410 ;
        RECT 52.055 34.910 52.225 35.410 ;
        RECT 55.055 35.120 57.215 35.470 ;
        RECT 68.055 35.120 70.215 35.470 ;
        RECT 48.425 34.680 48.885 34.850 ;
        RECT 21.805 34.190 23.965 34.540 ;
        RECT 34.805 34.190 36.965 34.540 ;
        RECT 55.055 34.290 57.215 34.640 ;
        RECT 68.055 34.290 70.215 34.640 ;
        RECT 21.805 33.360 23.965 33.710 ;
        RECT 34.805 33.360 36.965 33.710 ;
        RECT 55.055 33.460 57.215 33.810 ;
        RECT 68.055 33.460 70.215 33.810 ;
        RECT 21.805 32.530 23.965 32.880 ;
        RECT 34.805 32.530 36.965 32.880 ;
        RECT 40.325 32.240 40.495 32.740 ;
        RECT 41.385 32.240 41.555 32.740 ;
        RECT 43.715 32.240 43.885 32.740 ;
        RECT 44.775 32.240 44.945 32.740 ;
        RECT 48.425 32.690 48.885 32.860 ;
        RECT 51.425 32.690 51.885 32.860 ;
        RECT 55.055 32.630 57.215 32.980 ;
        RECT 68.055 32.630 70.215 32.980 ;
        RECT 21.805 31.700 23.965 32.050 ;
        RECT 34.805 31.700 36.965 32.050 ;
        RECT 40.710 32.010 41.170 32.180 ;
        RECT 44.100 32.010 44.560 32.180 ;
        RECT 48.085 32.130 48.255 32.630 ;
        RECT 49.055 32.130 49.225 32.630 ;
        RECT 51.085 32.130 51.255 32.630 ;
        RECT 52.055 32.130 52.225 32.630 ;
        RECT 48.425 31.900 48.885 32.070 ;
        RECT 55.055 31.800 57.215 32.150 ;
        RECT 68.055 31.800 70.215 32.150 ;
        RECT 21.805 30.870 23.965 31.220 ;
        RECT 34.805 30.870 36.965 31.220 ;
        RECT 55.055 30.970 57.215 31.320 ;
        RECT 68.055 30.970 70.215 31.320 ;
        RECT 21.805 30.040 23.965 30.390 ;
        RECT 34.805 30.040 36.965 30.390 ;
        RECT 55.055 30.140 57.215 30.490 ;
        RECT 68.055 30.140 70.215 30.490 ;
        RECT 48.435 29.910 48.895 30.080 ;
        RECT 51.425 29.910 51.885 30.080 ;
        RECT 21.805 29.210 23.965 29.560 ;
        RECT 34.805 29.210 36.965 29.560 ;
        RECT 48.095 29.350 48.265 29.850 ;
        RECT 49.065 29.350 49.235 29.850 ;
        RECT 51.085 29.350 51.255 29.850 ;
        RECT 52.055 29.350 52.225 29.850 ;
        RECT 55.055 29.310 57.215 29.660 ;
        RECT 68.055 29.310 70.215 29.660 ;
        RECT 48.435 29.120 48.895 29.290 ;
        RECT 21.805 28.380 23.965 28.730 ;
        RECT 34.805 28.380 36.965 28.730 ;
        RECT 55.055 28.480 57.215 28.830 ;
        RECT 68.055 28.480 70.215 28.830 ;
        RECT 21.805 27.550 23.965 27.900 ;
        RECT 34.805 27.550 36.965 27.900 ;
        RECT 55.055 27.650 57.215 28.000 ;
        RECT 68.055 27.650 70.215 28.000 ;
        RECT 48.435 27.130 48.895 27.300 ;
        RECT 21.805 26.720 23.965 27.070 ;
        RECT 34.805 26.720 36.965 27.070 ;
        RECT 48.095 26.570 48.265 27.070 ;
        RECT 49.065 26.570 49.235 27.070 ;
        RECT 55.055 26.820 57.215 27.170 ;
        RECT 68.055 26.820 70.215 27.170 ;
        RECT 21.805 25.890 23.965 26.240 ;
        RECT 34.805 25.890 36.965 26.240 ;
        RECT 55.055 25.990 57.215 26.340 ;
        RECT 68.055 25.990 70.215 26.340 ;
        RECT 21.805 25.060 23.965 25.410 ;
        RECT 34.805 25.060 36.965 25.410 ;
        RECT 55.055 25.160 57.215 25.510 ;
        RECT 68.055 25.160 70.215 25.510 ;
        RECT 21.805 24.230 23.965 24.580 ;
        RECT 34.805 24.230 36.965 24.580 ;
        RECT 55.055 24.330 57.215 24.680 ;
        RECT 68.055 24.330 70.215 24.680 ;
        RECT 21.805 23.400 23.965 23.750 ;
        RECT 34.805 23.400 36.965 23.750 ;
        RECT 55.055 23.500 57.215 23.850 ;
        RECT 68.055 23.500 70.215 23.850 ;
        RECT 21.805 22.570 23.965 22.920 ;
        RECT 34.805 22.570 36.965 22.920 ;
        RECT 68.055 22.670 70.215 23.020 ;
      LAYER mcon ;
        RECT 42.775 79.510 42.945 79.680 ;
        RECT 43.300 79.290 43.470 79.460 ;
        RECT 48.595 79.545 48.765 79.715 ;
        RECT 45.455 79.305 45.625 79.475 ;
        RECT 21.905 78.270 22.075 78.440 ;
        RECT 22.265 78.270 22.435 78.440 ;
        RECT 22.625 78.270 22.795 78.440 ;
        RECT 22.985 78.270 23.155 78.440 ;
        RECT 23.345 78.270 23.515 78.440 ;
        RECT 23.705 78.270 23.875 78.440 ;
        RECT 34.900 78.270 35.070 78.440 ;
        RECT 35.260 78.270 35.430 78.440 ;
        RECT 35.620 78.270 35.790 78.440 ;
        RECT 35.980 78.270 36.150 78.440 ;
        RECT 36.340 78.270 36.510 78.440 ;
        RECT 36.700 78.270 36.870 78.440 ;
        RECT 55.155 78.370 55.325 78.540 ;
        RECT 55.515 78.370 55.685 78.540 ;
        RECT 55.875 78.370 56.045 78.540 ;
        RECT 56.235 78.370 56.405 78.540 ;
        RECT 56.595 78.370 56.765 78.540 ;
        RECT 56.955 78.370 57.125 78.540 ;
        RECT 68.150 78.370 68.320 78.540 ;
        RECT 68.510 78.370 68.680 78.540 ;
        RECT 68.870 78.370 69.040 78.540 ;
        RECT 69.230 78.370 69.400 78.540 ;
        RECT 69.590 78.370 69.760 78.540 ;
        RECT 69.950 78.370 70.120 78.540 ;
        RECT 21.905 77.440 22.075 77.610 ;
        RECT 22.265 77.440 22.435 77.610 ;
        RECT 22.625 77.440 22.795 77.610 ;
        RECT 22.985 77.440 23.155 77.610 ;
        RECT 23.345 77.440 23.515 77.610 ;
        RECT 23.705 77.440 23.875 77.610 ;
        RECT 34.900 77.440 35.070 77.610 ;
        RECT 35.260 77.440 35.430 77.610 ;
        RECT 35.620 77.440 35.790 77.610 ;
        RECT 35.980 77.440 36.150 77.610 ;
        RECT 36.340 77.440 36.510 77.610 ;
        RECT 36.700 77.440 36.870 77.610 ;
        RECT 55.155 77.540 55.325 77.710 ;
        RECT 55.515 77.540 55.685 77.710 ;
        RECT 55.875 77.540 56.045 77.710 ;
        RECT 56.235 77.540 56.405 77.710 ;
        RECT 56.595 77.540 56.765 77.710 ;
        RECT 56.955 77.540 57.125 77.710 ;
        RECT 68.150 77.540 68.320 77.710 ;
        RECT 68.510 77.540 68.680 77.710 ;
        RECT 68.870 77.540 69.040 77.710 ;
        RECT 69.230 77.540 69.400 77.710 ;
        RECT 69.590 77.540 69.760 77.710 ;
        RECT 69.950 77.540 70.120 77.710 ;
        RECT 21.905 76.610 22.075 76.780 ;
        RECT 22.265 76.610 22.435 76.780 ;
        RECT 22.625 76.610 22.795 76.780 ;
        RECT 22.985 76.610 23.155 76.780 ;
        RECT 23.345 76.610 23.515 76.780 ;
        RECT 23.705 76.610 23.875 76.780 ;
        RECT 34.900 76.610 35.070 76.780 ;
        RECT 35.260 76.610 35.430 76.780 ;
        RECT 35.620 76.610 35.790 76.780 ;
        RECT 35.980 76.610 36.150 76.780 ;
        RECT 36.340 76.610 36.510 76.780 ;
        RECT 36.700 76.610 36.870 76.780 ;
        RECT 46.815 76.705 46.985 76.875 ;
        RECT 55.155 76.710 55.325 76.880 ;
        RECT 55.515 76.710 55.685 76.880 ;
        RECT 55.875 76.710 56.045 76.880 ;
        RECT 56.235 76.710 56.405 76.880 ;
        RECT 56.595 76.710 56.765 76.880 ;
        RECT 56.955 76.710 57.125 76.880 ;
        RECT 68.150 76.710 68.320 76.880 ;
        RECT 68.510 76.710 68.680 76.880 ;
        RECT 68.870 76.710 69.040 76.880 ;
        RECT 69.230 76.710 69.400 76.880 ;
        RECT 69.590 76.710 69.760 76.880 ;
        RECT 69.950 76.710 70.120 76.880 ;
        RECT 21.905 75.780 22.075 75.950 ;
        RECT 22.265 75.780 22.435 75.950 ;
        RECT 22.625 75.780 22.795 75.950 ;
        RECT 22.985 75.780 23.155 75.950 ;
        RECT 23.345 75.780 23.515 75.950 ;
        RECT 23.705 75.780 23.875 75.950 ;
        RECT 34.900 75.780 35.070 75.950 ;
        RECT 35.260 75.780 35.430 75.950 ;
        RECT 35.620 75.780 35.790 75.950 ;
        RECT 35.980 75.780 36.150 75.950 ;
        RECT 36.340 75.780 36.510 75.950 ;
        RECT 36.700 75.780 36.870 75.950 ;
        RECT 55.155 75.880 55.325 76.050 ;
        RECT 55.515 75.880 55.685 76.050 ;
        RECT 55.875 75.880 56.045 76.050 ;
        RECT 56.235 75.880 56.405 76.050 ;
        RECT 56.595 75.880 56.765 76.050 ;
        RECT 56.955 75.880 57.125 76.050 ;
        RECT 68.150 75.880 68.320 76.050 ;
        RECT 68.510 75.880 68.680 76.050 ;
        RECT 68.870 75.880 69.040 76.050 ;
        RECT 69.230 75.880 69.400 76.050 ;
        RECT 69.590 75.880 69.760 76.050 ;
        RECT 69.950 75.880 70.120 76.050 ;
        RECT 21.905 74.950 22.075 75.120 ;
        RECT 22.265 74.950 22.435 75.120 ;
        RECT 22.625 74.950 22.795 75.120 ;
        RECT 22.985 74.950 23.155 75.120 ;
        RECT 23.345 74.950 23.515 75.120 ;
        RECT 23.705 74.950 23.875 75.120 ;
        RECT 43.800 75.120 43.970 75.290 ;
        RECT 44.160 75.120 44.330 75.290 ;
        RECT 46.990 75.120 47.160 75.290 ;
        RECT 47.350 75.120 47.520 75.290 ;
        RECT 34.900 74.950 35.070 75.120 ;
        RECT 35.260 74.950 35.430 75.120 ;
        RECT 35.620 74.950 35.790 75.120 ;
        RECT 35.980 74.950 36.150 75.120 ;
        RECT 36.340 74.950 36.510 75.120 ;
        RECT 36.700 74.950 36.870 75.120 ;
        RECT 55.155 75.050 55.325 75.220 ;
        RECT 55.515 75.050 55.685 75.220 ;
        RECT 55.875 75.050 56.045 75.220 ;
        RECT 56.235 75.050 56.405 75.220 ;
        RECT 56.595 75.050 56.765 75.220 ;
        RECT 56.955 75.050 57.125 75.220 ;
        RECT 68.150 75.050 68.320 75.220 ;
        RECT 68.510 75.050 68.680 75.220 ;
        RECT 68.870 75.050 69.040 75.220 ;
        RECT 69.230 75.050 69.400 75.220 ;
        RECT 69.590 75.050 69.760 75.220 ;
        RECT 69.950 75.050 70.120 75.220 ;
        RECT 21.905 74.120 22.075 74.290 ;
        RECT 22.265 74.120 22.435 74.290 ;
        RECT 22.625 74.120 22.795 74.290 ;
        RECT 22.985 74.120 23.155 74.290 ;
        RECT 23.345 74.120 23.515 74.290 ;
        RECT 23.705 74.120 23.875 74.290 ;
        RECT 34.900 74.120 35.070 74.290 ;
        RECT 35.260 74.120 35.430 74.290 ;
        RECT 35.620 74.120 35.790 74.290 ;
        RECT 35.980 74.120 36.150 74.290 ;
        RECT 36.340 74.120 36.510 74.290 ;
        RECT 36.700 74.120 36.870 74.290 ;
        RECT 55.155 74.220 55.325 74.390 ;
        RECT 55.515 74.220 55.685 74.390 ;
        RECT 55.875 74.220 56.045 74.390 ;
        RECT 56.235 74.220 56.405 74.390 ;
        RECT 56.595 74.220 56.765 74.390 ;
        RECT 56.955 74.220 57.125 74.390 ;
        RECT 68.150 74.220 68.320 74.390 ;
        RECT 68.510 74.220 68.680 74.390 ;
        RECT 68.870 74.220 69.040 74.390 ;
        RECT 69.230 74.220 69.400 74.390 ;
        RECT 69.590 74.220 69.760 74.390 ;
        RECT 69.950 74.220 70.120 74.390 ;
        RECT 21.905 73.290 22.075 73.460 ;
        RECT 22.265 73.290 22.435 73.460 ;
        RECT 22.625 73.290 22.795 73.460 ;
        RECT 22.985 73.290 23.155 73.460 ;
        RECT 23.345 73.290 23.515 73.460 ;
        RECT 23.705 73.290 23.875 73.460 ;
        RECT 34.900 73.290 35.070 73.460 ;
        RECT 35.260 73.290 35.430 73.460 ;
        RECT 35.620 73.290 35.790 73.460 ;
        RECT 35.980 73.290 36.150 73.460 ;
        RECT 36.340 73.290 36.510 73.460 ;
        RECT 36.700 73.290 36.870 73.460 ;
        RECT 55.155 73.390 55.325 73.560 ;
        RECT 55.515 73.390 55.685 73.560 ;
        RECT 55.875 73.390 56.045 73.560 ;
        RECT 56.235 73.390 56.405 73.560 ;
        RECT 56.595 73.390 56.765 73.560 ;
        RECT 56.955 73.390 57.125 73.560 ;
        RECT 68.150 73.390 68.320 73.560 ;
        RECT 68.510 73.390 68.680 73.560 ;
        RECT 68.870 73.390 69.040 73.560 ;
        RECT 69.230 73.390 69.400 73.560 ;
        RECT 69.590 73.390 69.760 73.560 ;
        RECT 69.950 73.390 70.120 73.560 ;
        RECT 21.905 72.460 22.075 72.630 ;
        RECT 22.265 72.460 22.435 72.630 ;
        RECT 22.625 72.460 22.795 72.630 ;
        RECT 22.985 72.460 23.155 72.630 ;
        RECT 23.345 72.460 23.515 72.630 ;
        RECT 23.705 72.460 23.875 72.630 ;
        RECT 34.900 72.460 35.070 72.630 ;
        RECT 35.260 72.460 35.430 72.630 ;
        RECT 35.620 72.460 35.790 72.630 ;
        RECT 35.980 72.460 36.150 72.630 ;
        RECT 36.340 72.460 36.510 72.630 ;
        RECT 36.700 72.460 36.870 72.630 ;
        RECT 55.155 72.560 55.325 72.730 ;
        RECT 55.515 72.560 55.685 72.730 ;
        RECT 55.875 72.560 56.045 72.730 ;
        RECT 56.235 72.560 56.405 72.730 ;
        RECT 56.595 72.560 56.765 72.730 ;
        RECT 56.955 72.560 57.125 72.730 ;
        RECT 68.150 72.560 68.320 72.730 ;
        RECT 68.510 72.560 68.680 72.730 ;
        RECT 68.870 72.560 69.040 72.730 ;
        RECT 69.230 72.560 69.400 72.730 ;
        RECT 69.590 72.560 69.760 72.730 ;
        RECT 69.950 72.560 70.120 72.730 ;
        RECT 21.905 71.630 22.075 71.800 ;
        RECT 22.265 71.630 22.435 71.800 ;
        RECT 22.625 71.630 22.795 71.800 ;
        RECT 22.985 71.630 23.155 71.800 ;
        RECT 23.345 71.630 23.515 71.800 ;
        RECT 23.705 71.630 23.875 71.800 ;
        RECT 34.900 71.630 35.070 71.800 ;
        RECT 35.260 71.630 35.430 71.800 ;
        RECT 35.620 71.630 35.790 71.800 ;
        RECT 35.980 71.630 36.150 71.800 ;
        RECT 36.340 71.630 36.510 71.800 ;
        RECT 36.700 71.630 36.870 71.800 ;
        RECT 42.485 71.750 42.655 71.920 ;
        RECT 55.155 71.730 55.325 71.900 ;
        RECT 55.515 71.730 55.685 71.900 ;
        RECT 55.875 71.730 56.045 71.900 ;
        RECT 56.235 71.730 56.405 71.900 ;
        RECT 56.595 71.730 56.765 71.900 ;
        RECT 56.955 71.730 57.125 71.900 ;
        RECT 68.150 71.730 68.320 71.900 ;
        RECT 68.510 71.730 68.680 71.900 ;
        RECT 68.870 71.730 69.040 71.900 ;
        RECT 69.230 71.730 69.400 71.900 ;
        RECT 69.590 71.730 69.760 71.900 ;
        RECT 69.950 71.730 70.120 71.900 ;
        RECT 21.905 70.800 22.075 70.970 ;
        RECT 22.265 70.800 22.435 70.970 ;
        RECT 22.625 70.800 22.795 70.970 ;
        RECT 22.985 70.800 23.155 70.970 ;
        RECT 23.345 70.800 23.515 70.970 ;
        RECT 23.705 70.800 23.875 70.970 ;
        RECT 34.900 70.800 35.070 70.970 ;
        RECT 35.260 70.800 35.430 70.970 ;
        RECT 35.620 70.800 35.790 70.970 ;
        RECT 35.980 70.800 36.150 70.970 ;
        RECT 36.340 70.800 36.510 70.970 ;
        RECT 36.700 70.800 36.870 70.970 ;
        RECT 55.155 70.900 55.325 71.070 ;
        RECT 55.515 70.900 55.685 71.070 ;
        RECT 55.875 70.900 56.045 71.070 ;
        RECT 56.235 70.900 56.405 71.070 ;
        RECT 56.595 70.900 56.765 71.070 ;
        RECT 56.955 70.900 57.125 71.070 ;
        RECT 68.150 70.900 68.320 71.070 ;
        RECT 68.510 70.900 68.680 71.070 ;
        RECT 68.870 70.900 69.040 71.070 ;
        RECT 69.230 70.900 69.400 71.070 ;
        RECT 69.590 70.900 69.760 71.070 ;
        RECT 69.950 70.900 70.120 71.070 ;
        RECT 21.905 69.970 22.075 70.140 ;
        RECT 22.265 69.970 22.435 70.140 ;
        RECT 22.625 69.970 22.795 70.140 ;
        RECT 22.985 69.970 23.155 70.140 ;
        RECT 23.345 69.970 23.515 70.140 ;
        RECT 23.705 69.970 23.875 70.140 ;
        RECT 34.900 69.970 35.070 70.140 ;
        RECT 35.260 69.970 35.430 70.140 ;
        RECT 35.620 69.970 35.790 70.140 ;
        RECT 35.980 69.970 36.150 70.140 ;
        RECT 36.340 69.970 36.510 70.140 ;
        RECT 36.700 69.970 36.870 70.140 ;
        RECT 55.155 70.070 55.325 70.240 ;
        RECT 55.515 70.070 55.685 70.240 ;
        RECT 55.875 70.070 56.045 70.240 ;
        RECT 56.235 70.070 56.405 70.240 ;
        RECT 56.595 70.070 56.765 70.240 ;
        RECT 56.955 70.070 57.125 70.240 ;
        RECT 68.150 70.070 68.320 70.240 ;
        RECT 68.510 70.070 68.680 70.240 ;
        RECT 68.870 70.070 69.040 70.240 ;
        RECT 69.230 70.070 69.400 70.240 ;
        RECT 69.590 70.070 69.760 70.240 ;
        RECT 69.950 70.070 70.120 70.240 ;
        RECT 21.905 69.140 22.075 69.310 ;
        RECT 22.265 69.140 22.435 69.310 ;
        RECT 22.625 69.140 22.795 69.310 ;
        RECT 22.985 69.140 23.155 69.310 ;
        RECT 23.345 69.140 23.515 69.310 ;
        RECT 23.705 69.140 23.875 69.310 ;
        RECT 34.900 69.140 35.070 69.310 ;
        RECT 35.260 69.140 35.430 69.310 ;
        RECT 35.620 69.140 35.790 69.310 ;
        RECT 35.980 69.140 36.150 69.310 ;
        RECT 36.340 69.140 36.510 69.310 ;
        RECT 36.700 69.140 36.870 69.310 ;
        RECT 55.155 69.240 55.325 69.410 ;
        RECT 55.515 69.240 55.685 69.410 ;
        RECT 55.875 69.240 56.045 69.410 ;
        RECT 56.235 69.240 56.405 69.410 ;
        RECT 56.595 69.240 56.765 69.410 ;
        RECT 56.955 69.240 57.125 69.410 ;
        RECT 68.150 69.240 68.320 69.410 ;
        RECT 68.510 69.240 68.680 69.410 ;
        RECT 68.870 69.240 69.040 69.410 ;
        RECT 69.230 69.240 69.400 69.410 ;
        RECT 69.590 69.240 69.760 69.410 ;
        RECT 69.950 69.240 70.120 69.410 ;
        RECT 21.905 68.310 22.075 68.480 ;
        RECT 22.265 68.310 22.435 68.480 ;
        RECT 22.625 68.310 22.795 68.480 ;
        RECT 22.985 68.310 23.155 68.480 ;
        RECT 23.345 68.310 23.515 68.480 ;
        RECT 23.705 68.310 23.875 68.480 ;
        RECT 34.900 68.310 35.070 68.480 ;
        RECT 35.260 68.310 35.430 68.480 ;
        RECT 35.620 68.310 35.790 68.480 ;
        RECT 35.980 68.310 36.150 68.480 ;
        RECT 36.340 68.310 36.510 68.480 ;
        RECT 36.700 68.310 36.870 68.480 ;
        RECT 55.155 68.410 55.325 68.580 ;
        RECT 55.515 68.410 55.685 68.580 ;
        RECT 55.875 68.410 56.045 68.580 ;
        RECT 56.235 68.410 56.405 68.580 ;
        RECT 56.595 68.410 56.765 68.580 ;
        RECT 56.955 68.410 57.125 68.580 ;
        RECT 68.150 68.410 68.320 68.580 ;
        RECT 68.510 68.410 68.680 68.580 ;
        RECT 68.870 68.410 69.040 68.580 ;
        RECT 69.230 68.410 69.400 68.580 ;
        RECT 69.590 68.410 69.760 68.580 ;
        RECT 69.950 68.410 70.120 68.580 ;
        RECT 21.905 67.480 22.075 67.650 ;
        RECT 22.265 67.480 22.435 67.650 ;
        RECT 22.625 67.480 22.795 67.650 ;
        RECT 22.985 67.480 23.155 67.650 ;
        RECT 23.345 67.480 23.515 67.650 ;
        RECT 23.705 67.480 23.875 67.650 ;
        RECT 34.900 67.480 35.070 67.650 ;
        RECT 35.260 67.480 35.430 67.650 ;
        RECT 35.620 67.480 35.790 67.650 ;
        RECT 35.980 67.480 36.150 67.650 ;
        RECT 36.340 67.480 36.510 67.650 ;
        RECT 36.700 67.480 36.870 67.650 ;
        RECT 45.875 67.470 46.045 67.640 ;
        RECT 49.215 67.500 49.385 67.670 ;
        RECT 55.155 67.580 55.325 67.750 ;
        RECT 55.515 67.580 55.685 67.750 ;
        RECT 55.875 67.580 56.045 67.750 ;
        RECT 56.235 67.580 56.405 67.750 ;
        RECT 56.595 67.580 56.765 67.750 ;
        RECT 56.955 67.580 57.125 67.750 ;
        RECT 68.150 67.580 68.320 67.750 ;
        RECT 68.510 67.580 68.680 67.750 ;
        RECT 68.870 67.580 69.040 67.750 ;
        RECT 69.230 67.580 69.400 67.750 ;
        RECT 69.590 67.580 69.760 67.750 ;
        RECT 69.950 67.580 70.120 67.750 ;
        RECT 45.345 67.075 45.515 67.245 ;
        RECT 46.405 67.075 46.575 67.245 ;
        RECT 48.685 67.105 48.855 67.275 ;
        RECT 49.745 67.105 49.915 67.275 ;
        RECT 21.905 66.650 22.075 66.820 ;
        RECT 22.265 66.650 22.435 66.820 ;
        RECT 22.625 66.650 22.795 66.820 ;
        RECT 22.985 66.650 23.155 66.820 ;
        RECT 23.345 66.650 23.515 66.820 ;
        RECT 23.705 66.650 23.875 66.820 ;
        RECT 34.900 66.650 35.070 66.820 ;
        RECT 35.260 66.650 35.430 66.820 ;
        RECT 35.620 66.650 35.790 66.820 ;
        RECT 35.980 66.650 36.150 66.820 ;
        RECT 36.340 66.650 36.510 66.820 ;
        RECT 36.700 66.650 36.870 66.820 ;
        RECT 42.360 66.670 42.530 66.840 ;
        RECT 45.875 66.680 46.045 66.850 ;
        RECT 55.155 66.750 55.325 66.920 ;
        RECT 55.515 66.750 55.685 66.920 ;
        RECT 55.875 66.750 56.045 66.920 ;
        RECT 56.235 66.750 56.405 66.920 ;
        RECT 56.595 66.750 56.765 66.920 ;
        RECT 56.955 66.750 57.125 66.920 ;
        RECT 68.150 66.750 68.320 66.920 ;
        RECT 68.510 66.750 68.680 66.920 ;
        RECT 68.870 66.750 69.040 66.920 ;
        RECT 69.230 66.750 69.400 66.920 ;
        RECT 69.590 66.750 69.760 66.920 ;
        RECT 69.950 66.750 70.120 66.920 ;
        RECT 21.905 65.820 22.075 65.990 ;
        RECT 22.265 65.820 22.435 65.990 ;
        RECT 22.625 65.820 22.795 65.990 ;
        RECT 22.985 65.820 23.155 65.990 ;
        RECT 23.345 65.820 23.515 65.990 ;
        RECT 23.705 65.820 23.875 65.990 ;
        RECT 34.900 65.820 35.070 65.990 ;
        RECT 35.260 65.820 35.430 65.990 ;
        RECT 35.620 65.820 35.790 65.990 ;
        RECT 35.980 65.820 36.150 65.990 ;
        RECT 36.340 65.820 36.510 65.990 ;
        RECT 36.700 65.820 36.870 65.990 ;
        RECT 55.155 65.920 55.325 66.090 ;
        RECT 55.515 65.920 55.685 66.090 ;
        RECT 55.875 65.920 56.045 66.090 ;
        RECT 56.235 65.920 56.405 66.090 ;
        RECT 56.595 65.920 56.765 66.090 ;
        RECT 56.955 65.920 57.125 66.090 ;
        RECT 68.150 65.920 68.320 66.090 ;
        RECT 68.510 65.920 68.680 66.090 ;
        RECT 68.870 65.920 69.040 66.090 ;
        RECT 69.230 65.920 69.400 66.090 ;
        RECT 69.590 65.920 69.760 66.090 ;
        RECT 69.950 65.920 70.120 66.090 ;
        RECT 21.905 64.990 22.075 65.160 ;
        RECT 22.265 64.990 22.435 65.160 ;
        RECT 22.625 64.990 22.795 65.160 ;
        RECT 22.985 64.990 23.155 65.160 ;
        RECT 23.345 64.990 23.515 65.160 ;
        RECT 23.705 64.990 23.875 65.160 ;
        RECT 34.900 64.990 35.070 65.160 ;
        RECT 35.260 64.990 35.430 65.160 ;
        RECT 35.620 64.990 35.790 65.160 ;
        RECT 35.980 64.990 36.150 65.160 ;
        RECT 36.340 64.990 36.510 65.160 ;
        RECT 36.700 64.990 36.870 65.160 ;
        RECT 55.155 65.090 55.325 65.260 ;
        RECT 55.515 65.090 55.685 65.260 ;
        RECT 55.875 65.090 56.045 65.260 ;
        RECT 56.235 65.090 56.405 65.260 ;
        RECT 56.595 65.090 56.765 65.260 ;
        RECT 56.955 65.090 57.125 65.260 ;
        RECT 68.150 65.090 68.320 65.260 ;
        RECT 68.510 65.090 68.680 65.260 ;
        RECT 68.870 65.090 69.040 65.260 ;
        RECT 69.230 65.090 69.400 65.260 ;
        RECT 69.590 65.090 69.760 65.260 ;
        RECT 69.950 65.090 70.120 65.260 ;
        RECT 42.370 64.430 42.540 64.600 ;
        RECT 45.865 64.420 46.035 64.590 ;
        RECT 21.905 64.160 22.075 64.330 ;
        RECT 22.265 64.160 22.435 64.330 ;
        RECT 22.625 64.160 22.795 64.330 ;
        RECT 22.985 64.160 23.155 64.330 ;
        RECT 23.345 64.160 23.515 64.330 ;
        RECT 23.705 64.160 23.875 64.330 ;
        RECT 34.900 64.160 35.070 64.330 ;
        RECT 35.260 64.160 35.430 64.330 ;
        RECT 35.620 64.160 35.790 64.330 ;
        RECT 35.980 64.160 36.150 64.330 ;
        RECT 36.340 64.160 36.510 64.330 ;
        RECT 36.700 64.160 36.870 64.330 ;
        RECT 41.885 64.035 42.055 64.205 ;
        RECT 42.855 64.035 43.025 64.205 ;
        RECT 45.335 64.025 45.505 64.195 ;
        RECT 46.395 64.025 46.565 64.195 ;
        RECT 48.685 64.025 48.855 64.195 ;
        RECT 49.745 64.025 49.915 64.195 ;
        RECT 55.155 64.260 55.325 64.430 ;
        RECT 55.515 64.260 55.685 64.430 ;
        RECT 55.875 64.260 56.045 64.430 ;
        RECT 56.235 64.260 56.405 64.430 ;
        RECT 56.595 64.260 56.765 64.430 ;
        RECT 56.955 64.260 57.125 64.430 ;
        RECT 68.150 64.260 68.320 64.430 ;
        RECT 68.510 64.260 68.680 64.430 ;
        RECT 68.870 64.260 69.040 64.430 ;
        RECT 69.230 64.260 69.400 64.430 ;
        RECT 69.590 64.260 69.760 64.430 ;
        RECT 69.950 64.260 70.120 64.430 ;
        RECT 45.865 63.630 46.035 63.800 ;
        RECT 49.215 63.630 49.385 63.800 ;
        RECT 21.905 63.330 22.075 63.500 ;
        RECT 22.265 63.330 22.435 63.500 ;
        RECT 22.625 63.330 22.795 63.500 ;
        RECT 22.985 63.330 23.155 63.500 ;
        RECT 23.345 63.330 23.515 63.500 ;
        RECT 23.705 63.330 23.875 63.500 ;
        RECT 34.900 63.330 35.070 63.500 ;
        RECT 35.260 63.330 35.430 63.500 ;
        RECT 35.620 63.330 35.790 63.500 ;
        RECT 35.980 63.330 36.150 63.500 ;
        RECT 36.340 63.330 36.510 63.500 ;
        RECT 36.700 63.330 36.870 63.500 ;
        RECT 55.155 63.430 55.325 63.600 ;
        RECT 55.515 63.430 55.685 63.600 ;
        RECT 55.875 63.430 56.045 63.600 ;
        RECT 56.235 63.430 56.405 63.600 ;
        RECT 56.595 63.430 56.765 63.600 ;
        RECT 56.955 63.430 57.125 63.600 ;
        RECT 68.150 63.430 68.320 63.600 ;
        RECT 68.510 63.430 68.680 63.600 ;
        RECT 68.870 63.430 69.040 63.600 ;
        RECT 69.230 63.430 69.400 63.600 ;
        RECT 69.590 63.430 69.760 63.600 ;
        RECT 69.950 63.430 70.120 63.600 ;
        RECT 21.905 62.500 22.075 62.670 ;
        RECT 22.265 62.500 22.435 62.670 ;
        RECT 22.625 62.500 22.795 62.670 ;
        RECT 22.985 62.500 23.155 62.670 ;
        RECT 23.345 62.500 23.515 62.670 ;
        RECT 23.705 62.500 23.875 62.670 ;
        RECT 34.900 62.500 35.070 62.670 ;
        RECT 35.260 62.500 35.430 62.670 ;
        RECT 35.620 62.500 35.790 62.670 ;
        RECT 35.980 62.500 36.150 62.670 ;
        RECT 36.340 62.500 36.510 62.670 ;
        RECT 36.700 62.500 36.870 62.670 ;
        RECT 55.155 62.600 55.325 62.770 ;
        RECT 55.515 62.600 55.685 62.770 ;
        RECT 55.875 62.600 56.045 62.770 ;
        RECT 56.235 62.600 56.405 62.770 ;
        RECT 56.595 62.600 56.765 62.770 ;
        RECT 56.955 62.600 57.125 62.770 ;
        RECT 68.150 62.600 68.320 62.770 ;
        RECT 68.510 62.600 68.680 62.770 ;
        RECT 68.870 62.600 69.040 62.770 ;
        RECT 69.230 62.600 69.400 62.770 ;
        RECT 69.590 62.600 69.760 62.770 ;
        RECT 69.950 62.600 70.120 62.770 ;
        RECT 21.905 61.670 22.075 61.840 ;
        RECT 22.265 61.670 22.435 61.840 ;
        RECT 22.625 61.670 22.795 61.840 ;
        RECT 22.985 61.670 23.155 61.840 ;
        RECT 23.345 61.670 23.515 61.840 ;
        RECT 23.705 61.670 23.875 61.840 ;
        RECT 34.900 61.670 35.070 61.840 ;
        RECT 35.260 61.670 35.430 61.840 ;
        RECT 35.620 61.670 35.790 61.840 ;
        RECT 35.980 61.670 36.150 61.840 ;
        RECT 36.340 61.670 36.510 61.840 ;
        RECT 36.700 61.670 36.870 61.840 ;
        RECT 55.155 61.770 55.325 61.940 ;
        RECT 55.515 61.770 55.685 61.940 ;
        RECT 55.875 61.770 56.045 61.940 ;
        RECT 56.235 61.770 56.405 61.940 ;
        RECT 56.595 61.770 56.765 61.940 ;
        RECT 56.955 61.770 57.125 61.940 ;
        RECT 68.150 61.770 68.320 61.940 ;
        RECT 68.510 61.770 68.680 61.940 ;
        RECT 68.870 61.770 69.040 61.940 ;
        RECT 69.230 61.770 69.400 61.940 ;
        RECT 69.590 61.770 69.760 61.940 ;
        RECT 69.950 61.770 70.120 61.940 ;
        RECT 21.905 60.840 22.075 61.010 ;
        RECT 22.265 60.840 22.435 61.010 ;
        RECT 22.625 60.840 22.795 61.010 ;
        RECT 22.985 60.840 23.155 61.010 ;
        RECT 23.345 60.840 23.515 61.010 ;
        RECT 23.705 60.840 23.875 61.010 ;
        RECT 34.900 60.840 35.070 61.010 ;
        RECT 35.260 60.840 35.430 61.010 ;
        RECT 35.620 60.840 35.790 61.010 ;
        RECT 35.980 60.840 36.150 61.010 ;
        RECT 36.340 60.840 36.510 61.010 ;
        RECT 36.700 60.840 36.870 61.010 ;
        RECT 55.155 60.940 55.325 61.110 ;
        RECT 55.515 60.940 55.685 61.110 ;
        RECT 55.875 60.940 56.045 61.110 ;
        RECT 56.235 60.940 56.405 61.110 ;
        RECT 56.595 60.940 56.765 61.110 ;
        RECT 56.955 60.940 57.125 61.110 ;
        RECT 68.150 60.940 68.320 61.110 ;
        RECT 68.510 60.940 68.680 61.110 ;
        RECT 68.870 60.940 69.040 61.110 ;
        RECT 69.230 60.940 69.400 61.110 ;
        RECT 69.590 60.940 69.760 61.110 ;
        RECT 69.950 60.940 70.120 61.110 ;
        RECT 21.905 60.010 22.075 60.180 ;
        RECT 22.265 60.010 22.435 60.180 ;
        RECT 22.625 60.010 22.795 60.180 ;
        RECT 22.985 60.010 23.155 60.180 ;
        RECT 23.345 60.010 23.515 60.180 ;
        RECT 23.705 60.010 23.875 60.180 ;
        RECT 34.900 60.010 35.070 60.180 ;
        RECT 35.260 60.010 35.430 60.180 ;
        RECT 35.620 60.010 35.790 60.180 ;
        RECT 35.980 60.010 36.150 60.180 ;
        RECT 36.340 60.010 36.510 60.180 ;
        RECT 36.700 60.010 36.870 60.180 ;
        RECT 55.155 60.110 55.325 60.280 ;
        RECT 55.515 60.110 55.685 60.280 ;
        RECT 55.875 60.110 56.045 60.280 ;
        RECT 56.235 60.110 56.405 60.280 ;
        RECT 56.595 60.110 56.765 60.280 ;
        RECT 56.955 60.110 57.125 60.280 ;
        RECT 68.150 60.110 68.320 60.280 ;
        RECT 68.510 60.110 68.680 60.280 ;
        RECT 68.870 60.110 69.040 60.280 ;
        RECT 69.230 60.110 69.400 60.280 ;
        RECT 69.590 60.110 69.760 60.280 ;
        RECT 69.950 60.110 70.120 60.280 ;
        RECT 21.905 59.180 22.075 59.350 ;
        RECT 22.265 59.180 22.435 59.350 ;
        RECT 22.625 59.180 22.795 59.350 ;
        RECT 22.985 59.180 23.155 59.350 ;
        RECT 23.345 59.180 23.515 59.350 ;
        RECT 23.705 59.180 23.875 59.350 ;
        RECT 34.900 59.180 35.070 59.350 ;
        RECT 35.260 59.180 35.430 59.350 ;
        RECT 35.620 59.180 35.790 59.350 ;
        RECT 35.980 59.180 36.150 59.350 ;
        RECT 36.340 59.180 36.510 59.350 ;
        RECT 36.700 59.180 36.870 59.350 ;
        RECT 55.155 59.280 55.325 59.450 ;
        RECT 55.515 59.280 55.685 59.450 ;
        RECT 55.875 59.280 56.045 59.450 ;
        RECT 56.235 59.280 56.405 59.450 ;
        RECT 56.595 59.280 56.765 59.450 ;
        RECT 56.955 59.280 57.125 59.450 ;
        RECT 68.150 59.280 68.320 59.450 ;
        RECT 68.510 59.280 68.680 59.450 ;
        RECT 68.870 59.280 69.040 59.450 ;
        RECT 69.230 59.280 69.400 59.450 ;
        RECT 69.590 59.280 69.760 59.450 ;
        RECT 69.950 59.280 70.120 59.450 ;
        RECT 44.245 58.710 44.415 58.880 ;
        RECT 48.580 58.650 48.750 58.820 ;
        RECT 51.580 58.650 51.750 58.820 ;
        RECT 21.905 58.350 22.075 58.520 ;
        RECT 22.265 58.350 22.435 58.520 ;
        RECT 22.625 58.350 22.795 58.520 ;
        RECT 22.985 58.350 23.155 58.520 ;
        RECT 23.345 58.350 23.515 58.520 ;
        RECT 23.705 58.350 23.875 58.520 ;
        RECT 34.900 58.350 35.070 58.520 ;
        RECT 35.260 58.350 35.430 58.520 ;
        RECT 35.620 58.350 35.790 58.520 ;
        RECT 35.980 58.350 36.150 58.520 ;
        RECT 36.340 58.350 36.510 58.520 ;
        RECT 36.700 58.350 36.870 58.520 ;
        RECT 43.715 58.315 43.885 58.485 ;
        RECT 44.775 58.315 44.945 58.485 ;
        RECT 51.095 58.255 51.265 58.425 ;
        RECT 52.065 58.255 52.235 58.425 ;
        RECT 55.155 58.450 55.325 58.620 ;
        RECT 55.515 58.450 55.685 58.620 ;
        RECT 55.875 58.450 56.045 58.620 ;
        RECT 56.235 58.450 56.405 58.620 ;
        RECT 56.595 58.450 56.765 58.620 ;
        RECT 56.955 58.450 57.125 58.620 ;
        RECT 68.150 58.450 68.320 58.620 ;
        RECT 68.510 58.450 68.680 58.620 ;
        RECT 68.870 58.450 69.040 58.620 ;
        RECT 69.230 58.450 69.400 58.620 ;
        RECT 69.590 58.450 69.760 58.620 ;
        RECT 69.950 58.450 70.120 58.620 ;
        RECT 48.580 57.860 48.750 58.030 ;
        RECT 21.905 57.520 22.075 57.690 ;
        RECT 22.265 57.520 22.435 57.690 ;
        RECT 22.625 57.520 22.795 57.690 ;
        RECT 22.985 57.520 23.155 57.690 ;
        RECT 23.345 57.520 23.515 57.690 ;
        RECT 23.705 57.520 23.875 57.690 ;
        RECT 34.900 57.520 35.070 57.690 ;
        RECT 35.260 57.520 35.430 57.690 ;
        RECT 35.620 57.520 35.790 57.690 ;
        RECT 35.980 57.520 36.150 57.690 ;
        RECT 36.340 57.520 36.510 57.690 ;
        RECT 36.700 57.520 36.870 57.690 ;
        RECT 55.155 57.620 55.325 57.790 ;
        RECT 55.515 57.620 55.685 57.790 ;
        RECT 55.875 57.620 56.045 57.790 ;
        RECT 56.235 57.620 56.405 57.790 ;
        RECT 56.595 57.620 56.765 57.790 ;
        RECT 56.955 57.620 57.125 57.790 ;
        RECT 68.150 57.620 68.320 57.790 ;
        RECT 68.510 57.620 68.680 57.790 ;
        RECT 68.870 57.620 69.040 57.790 ;
        RECT 69.230 57.620 69.400 57.790 ;
        RECT 69.590 57.620 69.760 57.790 ;
        RECT 69.950 57.620 70.120 57.790 ;
        RECT 21.905 56.690 22.075 56.860 ;
        RECT 22.265 56.690 22.435 56.860 ;
        RECT 22.625 56.690 22.795 56.860 ;
        RECT 22.985 56.690 23.155 56.860 ;
        RECT 23.345 56.690 23.515 56.860 ;
        RECT 23.705 56.690 23.875 56.860 ;
        RECT 34.900 56.690 35.070 56.860 ;
        RECT 35.260 56.690 35.430 56.860 ;
        RECT 35.620 56.690 35.790 56.860 ;
        RECT 35.980 56.690 36.150 56.860 ;
        RECT 36.340 56.690 36.510 56.860 ;
        RECT 36.700 56.690 36.870 56.860 ;
        RECT 55.155 56.790 55.325 56.960 ;
        RECT 55.515 56.790 55.685 56.960 ;
        RECT 55.875 56.790 56.045 56.960 ;
        RECT 56.235 56.790 56.405 56.960 ;
        RECT 56.595 56.790 56.765 56.960 ;
        RECT 56.955 56.790 57.125 56.960 ;
        RECT 68.150 56.790 68.320 56.960 ;
        RECT 68.510 56.790 68.680 56.960 ;
        RECT 68.870 56.790 69.040 56.960 ;
        RECT 69.230 56.790 69.400 56.960 ;
        RECT 69.590 56.790 69.760 56.960 ;
        RECT 69.950 56.790 70.120 56.960 ;
        RECT 21.905 55.860 22.075 56.030 ;
        RECT 22.265 55.860 22.435 56.030 ;
        RECT 22.625 55.860 22.795 56.030 ;
        RECT 22.985 55.860 23.155 56.030 ;
        RECT 23.345 55.860 23.515 56.030 ;
        RECT 23.705 55.860 23.875 56.030 ;
        RECT 34.900 55.860 35.070 56.030 ;
        RECT 35.260 55.860 35.430 56.030 ;
        RECT 35.620 55.860 35.790 56.030 ;
        RECT 35.980 55.860 36.150 56.030 ;
        RECT 36.340 55.860 36.510 56.030 ;
        RECT 36.700 55.860 36.870 56.030 ;
        RECT 55.155 55.960 55.325 56.130 ;
        RECT 55.515 55.960 55.685 56.130 ;
        RECT 55.875 55.960 56.045 56.130 ;
        RECT 56.235 55.960 56.405 56.130 ;
        RECT 56.595 55.960 56.765 56.130 ;
        RECT 56.955 55.960 57.125 56.130 ;
        RECT 68.150 55.960 68.320 56.130 ;
        RECT 68.510 55.960 68.680 56.130 ;
        RECT 68.870 55.960 69.040 56.130 ;
        RECT 69.230 55.960 69.400 56.130 ;
        RECT 69.590 55.960 69.760 56.130 ;
        RECT 69.950 55.960 70.120 56.130 ;
        RECT 21.905 55.030 22.075 55.200 ;
        RECT 22.265 55.030 22.435 55.200 ;
        RECT 22.625 55.030 22.795 55.200 ;
        RECT 22.985 55.030 23.155 55.200 ;
        RECT 23.345 55.030 23.515 55.200 ;
        RECT 23.705 55.030 23.875 55.200 ;
        RECT 34.900 55.030 35.070 55.200 ;
        RECT 35.260 55.030 35.430 55.200 ;
        RECT 35.620 55.030 35.790 55.200 ;
        RECT 35.980 55.030 36.150 55.200 ;
        RECT 36.340 55.030 36.510 55.200 ;
        RECT 36.700 55.030 36.870 55.200 ;
        RECT 55.155 55.130 55.325 55.300 ;
        RECT 55.515 55.130 55.685 55.300 ;
        RECT 55.875 55.130 56.045 55.300 ;
        RECT 56.235 55.130 56.405 55.300 ;
        RECT 56.595 55.130 56.765 55.300 ;
        RECT 56.955 55.130 57.125 55.300 ;
        RECT 68.150 55.130 68.320 55.300 ;
        RECT 68.510 55.130 68.680 55.300 ;
        RECT 68.870 55.130 69.040 55.300 ;
        RECT 69.230 55.130 69.400 55.300 ;
        RECT 69.590 55.130 69.760 55.300 ;
        RECT 69.950 55.130 70.120 55.300 ;
        RECT 21.905 54.200 22.075 54.370 ;
        RECT 22.265 54.200 22.435 54.370 ;
        RECT 22.625 54.200 22.795 54.370 ;
        RECT 22.985 54.200 23.155 54.370 ;
        RECT 23.345 54.200 23.515 54.370 ;
        RECT 23.705 54.200 23.875 54.370 ;
        RECT 34.900 54.200 35.070 54.370 ;
        RECT 35.260 54.200 35.430 54.370 ;
        RECT 35.620 54.200 35.790 54.370 ;
        RECT 35.980 54.200 36.150 54.370 ;
        RECT 36.340 54.200 36.510 54.370 ;
        RECT 36.700 54.200 36.870 54.370 ;
        RECT 44.245 54.360 44.415 54.530 ;
        RECT 55.155 54.300 55.325 54.470 ;
        RECT 55.515 54.300 55.685 54.470 ;
        RECT 55.875 54.300 56.045 54.470 ;
        RECT 56.235 54.300 56.405 54.470 ;
        RECT 56.595 54.300 56.765 54.470 ;
        RECT 56.955 54.300 57.125 54.470 ;
        RECT 40.325 53.965 40.495 54.135 ;
        RECT 41.385 53.965 41.555 54.135 ;
        RECT 43.715 53.965 43.885 54.135 ;
        RECT 68.150 54.300 68.320 54.470 ;
        RECT 68.510 54.300 68.680 54.470 ;
        RECT 68.870 54.300 69.040 54.470 ;
        RECT 69.230 54.300 69.400 54.470 ;
        RECT 69.590 54.300 69.760 54.470 ;
        RECT 69.950 54.300 70.120 54.470 ;
        RECT 44.775 53.965 44.945 54.135 ;
        RECT 21.905 53.370 22.075 53.540 ;
        RECT 22.265 53.370 22.435 53.540 ;
        RECT 22.625 53.370 22.795 53.540 ;
        RECT 22.985 53.370 23.155 53.540 ;
        RECT 23.345 53.370 23.515 53.540 ;
        RECT 23.705 53.370 23.875 53.540 ;
        RECT 40.855 53.570 41.025 53.740 ;
        RECT 44.245 53.570 44.415 53.740 ;
        RECT 34.900 53.370 35.070 53.540 ;
        RECT 35.260 53.370 35.430 53.540 ;
        RECT 35.620 53.370 35.790 53.540 ;
        RECT 35.980 53.370 36.150 53.540 ;
        RECT 36.340 53.370 36.510 53.540 ;
        RECT 36.700 53.370 36.870 53.540 ;
        RECT 55.155 53.470 55.325 53.640 ;
        RECT 55.515 53.470 55.685 53.640 ;
        RECT 55.875 53.470 56.045 53.640 ;
        RECT 56.235 53.470 56.405 53.640 ;
        RECT 56.595 53.470 56.765 53.640 ;
        RECT 56.955 53.470 57.125 53.640 ;
        RECT 68.150 53.470 68.320 53.640 ;
        RECT 68.510 53.470 68.680 53.640 ;
        RECT 68.870 53.470 69.040 53.640 ;
        RECT 69.230 53.470 69.400 53.640 ;
        RECT 69.590 53.470 69.760 53.640 ;
        RECT 69.950 53.470 70.120 53.640 ;
        RECT 21.905 52.540 22.075 52.710 ;
        RECT 22.265 52.540 22.435 52.710 ;
        RECT 22.625 52.540 22.795 52.710 ;
        RECT 22.985 52.540 23.155 52.710 ;
        RECT 23.345 52.540 23.515 52.710 ;
        RECT 23.705 52.540 23.875 52.710 ;
        RECT 34.900 52.540 35.070 52.710 ;
        RECT 35.260 52.540 35.430 52.710 ;
        RECT 35.620 52.540 35.790 52.710 ;
        RECT 35.980 52.540 36.150 52.710 ;
        RECT 36.340 52.540 36.510 52.710 ;
        RECT 36.700 52.540 36.870 52.710 ;
        RECT 55.155 52.640 55.325 52.810 ;
        RECT 55.515 52.640 55.685 52.810 ;
        RECT 55.875 52.640 56.045 52.810 ;
        RECT 56.235 52.640 56.405 52.810 ;
        RECT 56.595 52.640 56.765 52.810 ;
        RECT 56.955 52.640 57.125 52.810 ;
        RECT 68.150 52.640 68.320 52.810 ;
        RECT 68.510 52.640 68.680 52.810 ;
        RECT 68.870 52.640 69.040 52.810 ;
        RECT 69.230 52.640 69.400 52.810 ;
        RECT 69.590 52.640 69.760 52.810 ;
        RECT 69.950 52.640 70.120 52.810 ;
        RECT 48.570 52.150 48.740 52.320 ;
        RECT 51.570 52.150 51.740 52.320 ;
        RECT 21.905 51.710 22.075 51.880 ;
        RECT 22.265 51.710 22.435 51.880 ;
        RECT 22.625 51.710 22.795 51.880 ;
        RECT 22.985 51.710 23.155 51.880 ;
        RECT 23.345 51.710 23.515 51.880 ;
        RECT 23.705 51.710 23.875 51.880 ;
        RECT 34.900 51.710 35.070 51.880 ;
        RECT 35.260 51.710 35.430 51.880 ;
        RECT 35.620 51.710 35.790 51.880 ;
        RECT 35.980 51.710 36.150 51.880 ;
        RECT 36.340 51.710 36.510 51.880 ;
        RECT 36.700 51.710 36.870 51.880 ;
        RECT 48.085 51.755 48.255 51.925 ;
        RECT 49.055 51.755 49.225 51.925 ;
        RECT 51.085 51.755 51.255 51.925 ;
        RECT 52.055 51.755 52.225 51.925 ;
        RECT 55.155 51.810 55.325 51.980 ;
        RECT 55.515 51.810 55.685 51.980 ;
        RECT 55.875 51.810 56.045 51.980 ;
        RECT 56.235 51.810 56.405 51.980 ;
        RECT 56.595 51.810 56.765 51.980 ;
        RECT 56.955 51.810 57.125 51.980 ;
        RECT 68.150 51.810 68.320 51.980 ;
        RECT 68.510 51.810 68.680 51.980 ;
        RECT 68.870 51.810 69.040 51.980 ;
        RECT 69.230 51.810 69.400 51.980 ;
        RECT 69.590 51.810 69.760 51.980 ;
        RECT 69.950 51.810 70.120 51.980 ;
        RECT 44.245 51.280 44.415 51.450 ;
        RECT 48.570 51.360 48.740 51.530 ;
        RECT 21.905 50.880 22.075 51.050 ;
        RECT 22.265 50.880 22.435 51.050 ;
        RECT 22.625 50.880 22.795 51.050 ;
        RECT 22.985 50.880 23.155 51.050 ;
        RECT 23.345 50.880 23.515 51.050 ;
        RECT 23.705 50.880 23.875 51.050 ;
        RECT 34.900 50.880 35.070 51.050 ;
        RECT 35.260 50.880 35.430 51.050 ;
        RECT 35.620 50.880 35.790 51.050 ;
        RECT 35.980 50.880 36.150 51.050 ;
        RECT 36.340 50.880 36.510 51.050 ;
        RECT 36.700 50.880 36.870 51.050 ;
        RECT 40.325 50.885 40.495 51.055 ;
        RECT 41.385 50.885 41.555 51.055 ;
        RECT 43.715 50.885 43.885 51.055 ;
        RECT 44.775 50.885 44.945 51.055 ;
        RECT 55.155 50.980 55.325 51.150 ;
        RECT 55.515 50.980 55.685 51.150 ;
        RECT 55.875 50.980 56.045 51.150 ;
        RECT 56.235 50.980 56.405 51.150 ;
        RECT 56.595 50.980 56.765 51.150 ;
        RECT 56.955 50.980 57.125 51.150 ;
        RECT 68.150 50.980 68.320 51.150 ;
        RECT 68.510 50.980 68.680 51.150 ;
        RECT 68.870 50.980 69.040 51.150 ;
        RECT 69.230 50.980 69.400 51.150 ;
        RECT 69.590 50.980 69.760 51.150 ;
        RECT 69.950 50.980 70.120 51.150 ;
        RECT 40.855 50.490 41.025 50.660 ;
        RECT 44.245 50.490 44.415 50.660 ;
        RECT 21.905 50.050 22.075 50.220 ;
        RECT 22.265 50.050 22.435 50.220 ;
        RECT 22.625 50.050 22.795 50.220 ;
        RECT 22.985 50.050 23.155 50.220 ;
        RECT 23.345 50.050 23.515 50.220 ;
        RECT 23.705 50.050 23.875 50.220 ;
        RECT 34.900 50.050 35.070 50.220 ;
        RECT 35.260 50.050 35.430 50.220 ;
        RECT 35.620 50.050 35.790 50.220 ;
        RECT 35.980 50.050 36.150 50.220 ;
        RECT 36.340 50.050 36.510 50.220 ;
        RECT 36.700 50.050 36.870 50.220 ;
        RECT 55.155 50.150 55.325 50.320 ;
        RECT 55.515 50.150 55.685 50.320 ;
        RECT 55.875 50.150 56.045 50.320 ;
        RECT 56.235 50.150 56.405 50.320 ;
        RECT 56.595 50.150 56.765 50.320 ;
        RECT 56.955 50.150 57.125 50.320 ;
        RECT 68.150 50.150 68.320 50.320 ;
        RECT 68.510 50.150 68.680 50.320 ;
        RECT 68.870 50.150 69.040 50.320 ;
        RECT 69.230 50.150 69.400 50.320 ;
        RECT 69.590 50.150 69.760 50.320 ;
        RECT 69.950 50.150 70.120 50.320 ;
        RECT 21.905 49.220 22.075 49.390 ;
        RECT 22.265 49.220 22.435 49.390 ;
        RECT 22.625 49.220 22.795 49.390 ;
        RECT 22.985 49.220 23.155 49.390 ;
        RECT 23.345 49.220 23.515 49.390 ;
        RECT 23.705 49.220 23.875 49.390 ;
        RECT 34.900 49.220 35.070 49.390 ;
        RECT 35.260 49.220 35.430 49.390 ;
        RECT 35.620 49.220 35.790 49.390 ;
        RECT 35.980 49.220 36.150 49.390 ;
        RECT 36.340 49.220 36.510 49.390 ;
        RECT 36.700 49.220 36.870 49.390 ;
        RECT 48.570 49.370 48.740 49.540 ;
        RECT 51.570 49.370 51.740 49.540 ;
        RECT 55.155 49.320 55.325 49.490 ;
        RECT 55.515 49.320 55.685 49.490 ;
        RECT 55.875 49.320 56.045 49.490 ;
        RECT 56.235 49.320 56.405 49.490 ;
        RECT 56.595 49.320 56.765 49.490 ;
        RECT 56.955 49.320 57.125 49.490 ;
        RECT 48.085 48.975 48.255 49.145 ;
        RECT 49.055 48.975 49.225 49.145 ;
        RECT 51.085 48.975 51.255 49.145 ;
        RECT 68.150 49.320 68.320 49.490 ;
        RECT 68.510 49.320 68.680 49.490 ;
        RECT 68.870 49.320 69.040 49.490 ;
        RECT 69.230 49.320 69.400 49.490 ;
        RECT 69.590 49.320 69.760 49.490 ;
        RECT 69.950 49.320 70.120 49.490 ;
        RECT 52.055 48.975 52.225 49.145 ;
        RECT 21.905 48.390 22.075 48.560 ;
        RECT 22.265 48.390 22.435 48.560 ;
        RECT 22.625 48.390 22.795 48.560 ;
        RECT 22.985 48.390 23.155 48.560 ;
        RECT 23.345 48.390 23.515 48.560 ;
        RECT 23.705 48.390 23.875 48.560 ;
        RECT 48.570 48.580 48.740 48.750 ;
        RECT 34.900 48.390 35.070 48.560 ;
        RECT 35.260 48.390 35.430 48.560 ;
        RECT 35.620 48.390 35.790 48.560 ;
        RECT 35.980 48.390 36.150 48.560 ;
        RECT 36.340 48.390 36.510 48.560 ;
        RECT 36.700 48.390 36.870 48.560 ;
        RECT 55.155 48.490 55.325 48.660 ;
        RECT 55.515 48.490 55.685 48.660 ;
        RECT 55.875 48.490 56.045 48.660 ;
        RECT 56.235 48.490 56.405 48.660 ;
        RECT 56.595 48.490 56.765 48.660 ;
        RECT 56.955 48.490 57.125 48.660 ;
        RECT 68.150 48.490 68.320 48.660 ;
        RECT 68.510 48.490 68.680 48.660 ;
        RECT 68.870 48.490 69.040 48.660 ;
        RECT 69.230 48.490 69.400 48.660 ;
        RECT 69.590 48.490 69.760 48.660 ;
        RECT 69.950 48.490 70.120 48.660 ;
        RECT 44.245 48.200 44.415 48.370 ;
        RECT 21.905 47.560 22.075 47.730 ;
        RECT 22.265 47.560 22.435 47.730 ;
        RECT 22.625 47.560 22.795 47.730 ;
        RECT 22.985 47.560 23.155 47.730 ;
        RECT 23.345 47.560 23.515 47.730 ;
        RECT 23.705 47.560 23.875 47.730 ;
        RECT 34.900 47.560 35.070 47.730 ;
        RECT 35.260 47.560 35.430 47.730 ;
        RECT 35.620 47.560 35.790 47.730 ;
        RECT 35.980 47.560 36.150 47.730 ;
        RECT 36.340 47.560 36.510 47.730 ;
        RECT 36.700 47.560 36.870 47.730 ;
        RECT 40.325 47.805 40.495 47.975 ;
        RECT 41.385 47.805 41.555 47.975 ;
        RECT 43.715 47.805 43.885 47.975 ;
        RECT 44.775 47.805 44.945 47.975 ;
        RECT 55.155 47.660 55.325 47.830 ;
        RECT 55.515 47.660 55.685 47.830 ;
        RECT 55.875 47.660 56.045 47.830 ;
        RECT 56.235 47.660 56.405 47.830 ;
        RECT 56.595 47.660 56.765 47.830 ;
        RECT 56.955 47.660 57.125 47.830 ;
        RECT 40.855 47.410 41.025 47.580 ;
        RECT 44.245 47.410 44.415 47.580 ;
        RECT 68.150 47.660 68.320 47.830 ;
        RECT 68.510 47.660 68.680 47.830 ;
        RECT 68.870 47.660 69.040 47.830 ;
        RECT 69.230 47.660 69.400 47.830 ;
        RECT 69.590 47.660 69.760 47.830 ;
        RECT 69.950 47.660 70.120 47.830 ;
        RECT 21.905 46.730 22.075 46.900 ;
        RECT 22.265 46.730 22.435 46.900 ;
        RECT 22.625 46.730 22.795 46.900 ;
        RECT 22.985 46.730 23.155 46.900 ;
        RECT 23.345 46.730 23.515 46.900 ;
        RECT 23.705 46.730 23.875 46.900 ;
        RECT 34.900 46.730 35.070 46.900 ;
        RECT 35.260 46.730 35.430 46.900 ;
        RECT 35.620 46.730 35.790 46.900 ;
        RECT 35.980 46.730 36.150 46.900 ;
        RECT 36.340 46.730 36.510 46.900 ;
        RECT 36.700 46.730 36.870 46.900 ;
        RECT 55.155 46.830 55.325 47.000 ;
        RECT 55.515 46.830 55.685 47.000 ;
        RECT 55.875 46.830 56.045 47.000 ;
        RECT 56.235 46.830 56.405 47.000 ;
        RECT 56.595 46.830 56.765 47.000 ;
        RECT 56.955 46.830 57.125 47.000 ;
        RECT 48.570 46.590 48.740 46.760 ;
        RECT 51.570 46.590 51.740 46.760 ;
        RECT 68.150 46.830 68.320 47.000 ;
        RECT 68.510 46.830 68.680 47.000 ;
        RECT 68.870 46.830 69.040 47.000 ;
        RECT 69.230 46.830 69.400 47.000 ;
        RECT 69.590 46.830 69.760 47.000 ;
        RECT 69.950 46.830 70.120 47.000 ;
        RECT 48.085 46.195 48.255 46.365 ;
        RECT 21.905 45.900 22.075 46.070 ;
        RECT 22.265 45.900 22.435 46.070 ;
        RECT 22.625 45.900 22.795 46.070 ;
        RECT 22.985 45.900 23.155 46.070 ;
        RECT 23.345 45.900 23.515 46.070 ;
        RECT 23.705 45.900 23.875 46.070 ;
        RECT 34.900 45.900 35.070 46.070 ;
        RECT 35.260 45.900 35.430 46.070 ;
        RECT 35.620 45.900 35.790 46.070 ;
        RECT 35.980 45.900 36.150 46.070 ;
        RECT 36.340 45.900 36.510 46.070 ;
        RECT 36.700 45.900 36.870 46.070 ;
        RECT 49.055 46.195 49.225 46.365 ;
        RECT 51.085 46.195 51.255 46.365 ;
        RECT 52.055 46.195 52.225 46.365 ;
        RECT 55.155 46.000 55.325 46.170 ;
        RECT 55.515 46.000 55.685 46.170 ;
        RECT 55.875 46.000 56.045 46.170 ;
        RECT 56.235 46.000 56.405 46.170 ;
        RECT 56.595 46.000 56.765 46.170 ;
        RECT 56.955 46.000 57.125 46.170 ;
        RECT 48.570 45.800 48.740 45.970 ;
        RECT 68.150 46.000 68.320 46.170 ;
        RECT 68.510 46.000 68.680 46.170 ;
        RECT 68.870 46.000 69.040 46.170 ;
        RECT 69.230 46.000 69.400 46.170 ;
        RECT 69.590 46.000 69.760 46.170 ;
        RECT 69.950 46.000 70.120 46.170 ;
        RECT 21.905 45.070 22.075 45.240 ;
        RECT 22.265 45.070 22.435 45.240 ;
        RECT 22.625 45.070 22.795 45.240 ;
        RECT 22.985 45.070 23.155 45.240 ;
        RECT 23.345 45.070 23.515 45.240 ;
        RECT 23.705 45.070 23.875 45.240 ;
        RECT 34.900 45.070 35.070 45.240 ;
        RECT 35.260 45.070 35.430 45.240 ;
        RECT 35.620 45.070 35.790 45.240 ;
        RECT 35.980 45.070 36.150 45.240 ;
        RECT 36.340 45.070 36.510 45.240 ;
        RECT 36.700 45.070 36.870 45.240 ;
        RECT 44.245 45.120 44.415 45.290 ;
        RECT 55.155 45.170 55.325 45.340 ;
        RECT 55.515 45.170 55.685 45.340 ;
        RECT 55.875 45.170 56.045 45.340 ;
        RECT 56.235 45.170 56.405 45.340 ;
        RECT 56.595 45.170 56.765 45.340 ;
        RECT 56.955 45.170 57.125 45.340 ;
        RECT 68.150 45.170 68.320 45.340 ;
        RECT 68.510 45.170 68.680 45.340 ;
        RECT 68.870 45.170 69.040 45.340 ;
        RECT 69.230 45.170 69.400 45.340 ;
        RECT 69.590 45.170 69.760 45.340 ;
        RECT 69.950 45.170 70.120 45.340 ;
        RECT 40.325 44.725 40.495 44.895 ;
        RECT 41.385 44.725 41.555 44.895 ;
        RECT 43.715 44.725 43.885 44.895 ;
        RECT 44.775 44.725 44.945 44.895 ;
        RECT 21.905 44.240 22.075 44.410 ;
        RECT 22.265 44.240 22.435 44.410 ;
        RECT 22.625 44.240 22.795 44.410 ;
        RECT 22.985 44.240 23.155 44.410 ;
        RECT 23.345 44.240 23.515 44.410 ;
        RECT 23.705 44.240 23.875 44.410 ;
        RECT 34.900 44.240 35.070 44.410 ;
        RECT 35.260 44.240 35.430 44.410 ;
        RECT 35.620 44.240 35.790 44.410 ;
        RECT 35.980 44.240 36.150 44.410 ;
        RECT 36.340 44.240 36.510 44.410 ;
        RECT 36.700 44.240 36.870 44.410 ;
        RECT 40.855 44.330 41.025 44.500 ;
        RECT 44.245 44.330 44.415 44.500 ;
        RECT 55.155 44.340 55.325 44.510 ;
        RECT 55.515 44.340 55.685 44.510 ;
        RECT 55.875 44.340 56.045 44.510 ;
        RECT 56.235 44.340 56.405 44.510 ;
        RECT 56.595 44.340 56.765 44.510 ;
        RECT 56.955 44.340 57.125 44.510 ;
        RECT 68.150 44.340 68.320 44.510 ;
        RECT 68.510 44.340 68.680 44.510 ;
        RECT 68.870 44.340 69.040 44.510 ;
        RECT 69.230 44.340 69.400 44.510 ;
        RECT 69.590 44.340 69.760 44.510 ;
        RECT 69.950 44.340 70.120 44.510 ;
        RECT 48.570 43.810 48.740 43.980 ;
        RECT 51.570 43.810 51.740 43.980 ;
        RECT 21.905 43.410 22.075 43.580 ;
        RECT 22.265 43.410 22.435 43.580 ;
        RECT 22.625 43.410 22.795 43.580 ;
        RECT 22.985 43.410 23.155 43.580 ;
        RECT 23.345 43.410 23.515 43.580 ;
        RECT 23.705 43.410 23.875 43.580 ;
        RECT 34.900 43.410 35.070 43.580 ;
        RECT 35.260 43.410 35.430 43.580 ;
        RECT 35.620 43.410 35.790 43.580 ;
        RECT 35.980 43.410 36.150 43.580 ;
        RECT 36.340 43.410 36.510 43.580 ;
        RECT 36.700 43.410 36.870 43.580 ;
        RECT 48.085 43.415 48.255 43.585 ;
        RECT 49.055 43.415 49.225 43.585 ;
        RECT 51.085 43.415 51.255 43.585 ;
        RECT 52.055 43.415 52.225 43.585 ;
        RECT 55.155 43.510 55.325 43.680 ;
        RECT 55.515 43.510 55.685 43.680 ;
        RECT 55.875 43.510 56.045 43.680 ;
        RECT 56.235 43.510 56.405 43.680 ;
        RECT 56.595 43.510 56.765 43.680 ;
        RECT 56.955 43.510 57.125 43.680 ;
        RECT 68.150 43.510 68.320 43.680 ;
        RECT 68.510 43.510 68.680 43.680 ;
        RECT 68.870 43.510 69.040 43.680 ;
        RECT 69.230 43.510 69.400 43.680 ;
        RECT 69.590 43.510 69.760 43.680 ;
        RECT 69.950 43.510 70.120 43.680 ;
        RECT 48.570 43.020 48.740 43.190 ;
        RECT 21.905 42.580 22.075 42.750 ;
        RECT 22.265 42.580 22.435 42.750 ;
        RECT 22.625 42.580 22.795 42.750 ;
        RECT 22.985 42.580 23.155 42.750 ;
        RECT 23.345 42.580 23.515 42.750 ;
        RECT 23.705 42.580 23.875 42.750 ;
        RECT 34.900 42.580 35.070 42.750 ;
        RECT 35.260 42.580 35.430 42.750 ;
        RECT 35.620 42.580 35.790 42.750 ;
        RECT 35.980 42.580 36.150 42.750 ;
        RECT 36.340 42.580 36.510 42.750 ;
        RECT 36.700 42.580 36.870 42.750 ;
        RECT 55.155 42.680 55.325 42.850 ;
        RECT 55.515 42.680 55.685 42.850 ;
        RECT 55.875 42.680 56.045 42.850 ;
        RECT 56.235 42.680 56.405 42.850 ;
        RECT 56.595 42.680 56.765 42.850 ;
        RECT 56.955 42.680 57.125 42.850 ;
        RECT 68.150 42.680 68.320 42.850 ;
        RECT 68.510 42.680 68.680 42.850 ;
        RECT 68.870 42.680 69.040 42.850 ;
        RECT 69.230 42.680 69.400 42.850 ;
        RECT 69.590 42.680 69.760 42.850 ;
        RECT 69.950 42.680 70.120 42.850 ;
        RECT 44.245 42.040 44.415 42.210 ;
        RECT 21.905 41.750 22.075 41.920 ;
        RECT 22.265 41.750 22.435 41.920 ;
        RECT 22.625 41.750 22.795 41.920 ;
        RECT 22.985 41.750 23.155 41.920 ;
        RECT 23.345 41.750 23.515 41.920 ;
        RECT 23.705 41.750 23.875 41.920 ;
        RECT 34.900 41.750 35.070 41.920 ;
        RECT 35.260 41.750 35.430 41.920 ;
        RECT 35.620 41.750 35.790 41.920 ;
        RECT 35.980 41.750 36.150 41.920 ;
        RECT 36.340 41.750 36.510 41.920 ;
        RECT 36.700 41.750 36.870 41.920 ;
        RECT 40.325 41.645 40.495 41.815 ;
        RECT 41.385 41.645 41.555 41.815 ;
        RECT 43.715 41.645 43.885 41.815 ;
        RECT 44.775 41.645 44.945 41.815 ;
        RECT 55.155 41.850 55.325 42.020 ;
        RECT 55.515 41.850 55.685 42.020 ;
        RECT 55.875 41.850 56.045 42.020 ;
        RECT 56.235 41.850 56.405 42.020 ;
        RECT 56.595 41.850 56.765 42.020 ;
        RECT 56.955 41.850 57.125 42.020 ;
        RECT 68.150 41.850 68.320 42.020 ;
        RECT 68.510 41.850 68.680 42.020 ;
        RECT 68.870 41.850 69.040 42.020 ;
        RECT 69.230 41.850 69.400 42.020 ;
        RECT 69.590 41.850 69.760 42.020 ;
        RECT 69.950 41.850 70.120 42.020 ;
        RECT 40.855 41.250 41.025 41.420 ;
        RECT 44.245 41.250 44.415 41.420 ;
        RECT 21.905 40.920 22.075 41.090 ;
        RECT 22.265 40.920 22.435 41.090 ;
        RECT 22.625 40.920 22.795 41.090 ;
        RECT 22.985 40.920 23.155 41.090 ;
        RECT 23.345 40.920 23.515 41.090 ;
        RECT 23.705 40.920 23.875 41.090 ;
        RECT 34.900 40.920 35.070 41.090 ;
        RECT 35.260 40.920 35.430 41.090 ;
        RECT 35.620 40.920 35.790 41.090 ;
        RECT 35.980 40.920 36.150 41.090 ;
        RECT 36.340 40.920 36.510 41.090 ;
        RECT 36.700 40.920 36.870 41.090 ;
        RECT 48.570 41.030 48.740 41.200 ;
        RECT 51.570 41.030 51.740 41.200 ;
        RECT 55.155 41.020 55.325 41.190 ;
        RECT 55.515 41.020 55.685 41.190 ;
        RECT 55.875 41.020 56.045 41.190 ;
        RECT 56.235 41.020 56.405 41.190 ;
        RECT 56.595 41.020 56.765 41.190 ;
        RECT 56.955 41.020 57.125 41.190 ;
        RECT 48.085 40.635 48.255 40.805 ;
        RECT 49.055 40.635 49.225 40.805 ;
        RECT 51.085 40.635 51.255 40.805 ;
        RECT 68.150 41.020 68.320 41.190 ;
        RECT 68.510 41.020 68.680 41.190 ;
        RECT 68.870 41.020 69.040 41.190 ;
        RECT 69.230 41.020 69.400 41.190 ;
        RECT 69.590 41.020 69.760 41.190 ;
        RECT 69.950 41.020 70.120 41.190 ;
        RECT 52.055 40.635 52.225 40.805 ;
        RECT 21.905 40.090 22.075 40.260 ;
        RECT 22.265 40.090 22.435 40.260 ;
        RECT 22.625 40.090 22.795 40.260 ;
        RECT 22.985 40.090 23.155 40.260 ;
        RECT 23.345 40.090 23.515 40.260 ;
        RECT 23.705 40.090 23.875 40.260 ;
        RECT 34.900 40.090 35.070 40.260 ;
        RECT 35.260 40.090 35.430 40.260 ;
        RECT 35.620 40.090 35.790 40.260 ;
        RECT 35.980 40.090 36.150 40.260 ;
        RECT 36.340 40.090 36.510 40.260 ;
        RECT 36.700 40.090 36.870 40.260 ;
        RECT 48.570 40.240 48.740 40.410 ;
        RECT 55.155 40.190 55.325 40.360 ;
        RECT 55.515 40.190 55.685 40.360 ;
        RECT 55.875 40.190 56.045 40.360 ;
        RECT 56.235 40.190 56.405 40.360 ;
        RECT 56.595 40.190 56.765 40.360 ;
        RECT 56.955 40.190 57.125 40.360 ;
        RECT 68.150 40.190 68.320 40.360 ;
        RECT 68.510 40.190 68.680 40.360 ;
        RECT 68.870 40.190 69.040 40.360 ;
        RECT 69.230 40.190 69.400 40.360 ;
        RECT 69.590 40.190 69.760 40.360 ;
        RECT 69.950 40.190 70.120 40.360 ;
        RECT 21.905 39.260 22.075 39.430 ;
        RECT 22.265 39.260 22.435 39.430 ;
        RECT 22.625 39.260 22.795 39.430 ;
        RECT 22.985 39.260 23.155 39.430 ;
        RECT 23.345 39.260 23.515 39.430 ;
        RECT 23.705 39.260 23.875 39.430 ;
        RECT 34.900 39.260 35.070 39.430 ;
        RECT 35.260 39.260 35.430 39.430 ;
        RECT 35.620 39.260 35.790 39.430 ;
        RECT 35.980 39.260 36.150 39.430 ;
        RECT 36.340 39.260 36.510 39.430 ;
        RECT 36.700 39.260 36.870 39.430 ;
        RECT 55.155 39.360 55.325 39.530 ;
        RECT 55.515 39.360 55.685 39.530 ;
        RECT 55.875 39.360 56.045 39.530 ;
        RECT 56.235 39.360 56.405 39.530 ;
        RECT 56.595 39.360 56.765 39.530 ;
        RECT 56.955 39.360 57.125 39.530 ;
        RECT 68.150 39.360 68.320 39.530 ;
        RECT 68.510 39.360 68.680 39.530 ;
        RECT 68.870 39.360 69.040 39.530 ;
        RECT 69.230 39.360 69.400 39.530 ;
        RECT 69.590 39.360 69.760 39.530 ;
        RECT 69.950 39.360 70.120 39.530 ;
        RECT 44.245 38.960 44.415 39.130 ;
        RECT 21.905 38.430 22.075 38.600 ;
        RECT 22.265 38.430 22.435 38.600 ;
        RECT 22.625 38.430 22.795 38.600 ;
        RECT 22.985 38.430 23.155 38.600 ;
        RECT 23.345 38.430 23.515 38.600 ;
        RECT 23.705 38.430 23.875 38.600 ;
        RECT 34.900 38.430 35.070 38.600 ;
        RECT 35.260 38.430 35.430 38.600 ;
        RECT 35.620 38.430 35.790 38.600 ;
        RECT 35.980 38.430 36.150 38.600 ;
        RECT 36.340 38.430 36.510 38.600 ;
        RECT 36.700 38.430 36.870 38.600 ;
        RECT 40.325 38.565 40.495 38.735 ;
        RECT 41.385 38.565 41.555 38.735 ;
        RECT 43.715 38.565 43.885 38.735 ;
        RECT 44.775 38.565 44.945 38.735 ;
        RECT 55.155 38.530 55.325 38.700 ;
        RECT 55.515 38.530 55.685 38.700 ;
        RECT 55.875 38.530 56.045 38.700 ;
        RECT 56.235 38.530 56.405 38.700 ;
        RECT 56.595 38.530 56.765 38.700 ;
        RECT 56.955 38.530 57.125 38.700 ;
        RECT 68.150 38.530 68.320 38.700 ;
        RECT 68.510 38.530 68.680 38.700 ;
        RECT 68.870 38.530 69.040 38.700 ;
        RECT 69.230 38.530 69.400 38.700 ;
        RECT 69.590 38.530 69.760 38.700 ;
        RECT 69.950 38.530 70.120 38.700 ;
        RECT 40.855 38.170 41.025 38.340 ;
        RECT 44.245 38.170 44.415 38.340 ;
        RECT 48.570 38.250 48.740 38.420 ;
        RECT 51.570 38.250 51.740 38.420 ;
        RECT 21.905 37.600 22.075 37.770 ;
        RECT 22.265 37.600 22.435 37.770 ;
        RECT 22.625 37.600 22.795 37.770 ;
        RECT 22.985 37.600 23.155 37.770 ;
        RECT 23.345 37.600 23.515 37.770 ;
        RECT 23.705 37.600 23.875 37.770 ;
        RECT 34.900 37.600 35.070 37.770 ;
        RECT 35.260 37.600 35.430 37.770 ;
        RECT 35.620 37.600 35.790 37.770 ;
        RECT 35.980 37.600 36.150 37.770 ;
        RECT 36.340 37.600 36.510 37.770 ;
        RECT 36.700 37.600 36.870 37.770 ;
        RECT 48.085 37.855 48.255 38.025 ;
        RECT 49.055 37.855 49.225 38.025 ;
        RECT 51.085 37.855 51.255 38.025 ;
        RECT 52.055 37.855 52.225 38.025 ;
        RECT 55.155 37.700 55.325 37.870 ;
        RECT 55.515 37.700 55.685 37.870 ;
        RECT 55.875 37.700 56.045 37.870 ;
        RECT 56.235 37.700 56.405 37.870 ;
        RECT 56.595 37.700 56.765 37.870 ;
        RECT 56.955 37.700 57.125 37.870 ;
        RECT 48.570 37.460 48.740 37.630 ;
        RECT 68.150 37.700 68.320 37.870 ;
        RECT 68.510 37.700 68.680 37.870 ;
        RECT 68.870 37.700 69.040 37.870 ;
        RECT 69.230 37.700 69.400 37.870 ;
        RECT 69.590 37.700 69.760 37.870 ;
        RECT 69.950 37.700 70.120 37.870 ;
        RECT 21.905 36.770 22.075 36.940 ;
        RECT 22.265 36.770 22.435 36.940 ;
        RECT 22.625 36.770 22.795 36.940 ;
        RECT 22.985 36.770 23.155 36.940 ;
        RECT 23.345 36.770 23.515 36.940 ;
        RECT 23.705 36.770 23.875 36.940 ;
        RECT 34.900 36.770 35.070 36.940 ;
        RECT 35.260 36.770 35.430 36.940 ;
        RECT 35.620 36.770 35.790 36.940 ;
        RECT 35.980 36.770 36.150 36.940 ;
        RECT 36.340 36.770 36.510 36.940 ;
        RECT 36.700 36.770 36.870 36.940 ;
        RECT 55.155 36.870 55.325 37.040 ;
        RECT 55.515 36.870 55.685 37.040 ;
        RECT 55.875 36.870 56.045 37.040 ;
        RECT 56.235 36.870 56.405 37.040 ;
        RECT 56.595 36.870 56.765 37.040 ;
        RECT 56.955 36.870 57.125 37.040 ;
        RECT 68.150 36.870 68.320 37.040 ;
        RECT 68.510 36.870 68.680 37.040 ;
        RECT 68.870 36.870 69.040 37.040 ;
        RECT 69.230 36.870 69.400 37.040 ;
        RECT 69.590 36.870 69.760 37.040 ;
        RECT 69.950 36.870 70.120 37.040 ;
        RECT 21.905 35.940 22.075 36.110 ;
        RECT 22.265 35.940 22.435 36.110 ;
        RECT 22.625 35.940 22.795 36.110 ;
        RECT 22.985 35.940 23.155 36.110 ;
        RECT 23.345 35.940 23.515 36.110 ;
        RECT 23.705 35.940 23.875 36.110 ;
        RECT 34.900 35.940 35.070 36.110 ;
        RECT 35.260 35.940 35.430 36.110 ;
        RECT 35.620 35.940 35.790 36.110 ;
        RECT 35.980 35.940 36.150 36.110 ;
        RECT 36.340 35.940 36.510 36.110 ;
        RECT 36.700 35.940 36.870 36.110 ;
        RECT 44.245 35.880 44.415 36.050 ;
        RECT 55.155 36.040 55.325 36.210 ;
        RECT 55.515 36.040 55.685 36.210 ;
        RECT 55.875 36.040 56.045 36.210 ;
        RECT 56.235 36.040 56.405 36.210 ;
        RECT 56.595 36.040 56.765 36.210 ;
        RECT 56.955 36.040 57.125 36.210 ;
        RECT 68.150 36.040 68.320 36.210 ;
        RECT 68.510 36.040 68.680 36.210 ;
        RECT 68.870 36.040 69.040 36.210 ;
        RECT 69.230 36.040 69.400 36.210 ;
        RECT 69.590 36.040 69.760 36.210 ;
        RECT 69.950 36.040 70.120 36.210 ;
        RECT 40.325 35.485 40.495 35.655 ;
        RECT 21.905 35.110 22.075 35.280 ;
        RECT 22.265 35.110 22.435 35.280 ;
        RECT 22.625 35.110 22.795 35.280 ;
        RECT 22.985 35.110 23.155 35.280 ;
        RECT 23.345 35.110 23.515 35.280 ;
        RECT 23.705 35.110 23.875 35.280 ;
        RECT 41.385 35.485 41.555 35.655 ;
        RECT 43.715 35.485 43.885 35.655 ;
        RECT 44.775 35.485 44.945 35.655 ;
        RECT 48.570 35.470 48.740 35.640 ;
        RECT 51.570 35.470 51.740 35.640 ;
        RECT 34.900 35.110 35.070 35.280 ;
        RECT 35.260 35.110 35.430 35.280 ;
        RECT 35.620 35.110 35.790 35.280 ;
        RECT 35.980 35.110 36.150 35.280 ;
        RECT 36.340 35.110 36.510 35.280 ;
        RECT 36.700 35.110 36.870 35.280 ;
        RECT 40.855 35.090 41.025 35.260 ;
        RECT 44.245 35.090 44.415 35.260 ;
        RECT 48.085 35.075 48.255 35.245 ;
        RECT 49.055 35.075 49.225 35.245 ;
        RECT 51.085 35.075 51.255 35.245 ;
        RECT 52.055 35.075 52.225 35.245 ;
        RECT 55.155 35.210 55.325 35.380 ;
        RECT 55.515 35.210 55.685 35.380 ;
        RECT 55.875 35.210 56.045 35.380 ;
        RECT 56.235 35.210 56.405 35.380 ;
        RECT 56.595 35.210 56.765 35.380 ;
        RECT 56.955 35.210 57.125 35.380 ;
        RECT 68.150 35.210 68.320 35.380 ;
        RECT 68.510 35.210 68.680 35.380 ;
        RECT 68.870 35.210 69.040 35.380 ;
        RECT 69.230 35.210 69.400 35.380 ;
        RECT 69.590 35.210 69.760 35.380 ;
        RECT 69.950 35.210 70.120 35.380 ;
        RECT 48.570 34.680 48.740 34.850 ;
        RECT 21.905 34.280 22.075 34.450 ;
        RECT 22.265 34.280 22.435 34.450 ;
        RECT 22.625 34.280 22.795 34.450 ;
        RECT 22.985 34.280 23.155 34.450 ;
        RECT 23.345 34.280 23.515 34.450 ;
        RECT 23.705 34.280 23.875 34.450 ;
        RECT 34.900 34.280 35.070 34.450 ;
        RECT 35.260 34.280 35.430 34.450 ;
        RECT 35.620 34.280 35.790 34.450 ;
        RECT 35.980 34.280 36.150 34.450 ;
        RECT 36.340 34.280 36.510 34.450 ;
        RECT 36.700 34.280 36.870 34.450 ;
        RECT 55.155 34.380 55.325 34.550 ;
        RECT 55.515 34.380 55.685 34.550 ;
        RECT 55.875 34.380 56.045 34.550 ;
        RECT 56.235 34.380 56.405 34.550 ;
        RECT 56.595 34.380 56.765 34.550 ;
        RECT 56.955 34.380 57.125 34.550 ;
        RECT 68.150 34.380 68.320 34.550 ;
        RECT 68.510 34.380 68.680 34.550 ;
        RECT 68.870 34.380 69.040 34.550 ;
        RECT 69.230 34.380 69.400 34.550 ;
        RECT 69.590 34.380 69.760 34.550 ;
        RECT 69.950 34.380 70.120 34.550 ;
        RECT 21.905 33.450 22.075 33.620 ;
        RECT 22.265 33.450 22.435 33.620 ;
        RECT 22.625 33.450 22.795 33.620 ;
        RECT 22.985 33.450 23.155 33.620 ;
        RECT 23.345 33.450 23.515 33.620 ;
        RECT 23.705 33.450 23.875 33.620 ;
        RECT 34.900 33.450 35.070 33.620 ;
        RECT 35.260 33.450 35.430 33.620 ;
        RECT 35.620 33.450 35.790 33.620 ;
        RECT 35.980 33.450 36.150 33.620 ;
        RECT 36.340 33.450 36.510 33.620 ;
        RECT 36.700 33.450 36.870 33.620 ;
        RECT 55.155 33.550 55.325 33.720 ;
        RECT 55.515 33.550 55.685 33.720 ;
        RECT 55.875 33.550 56.045 33.720 ;
        RECT 56.235 33.550 56.405 33.720 ;
        RECT 56.595 33.550 56.765 33.720 ;
        RECT 56.955 33.550 57.125 33.720 ;
        RECT 68.150 33.550 68.320 33.720 ;
        RECT 68.510 33.550 68.680 33.720 ;
        RECT 68.870 33.550 69.040 33.720 ;
        RECT 69.230 33.550 69.400 33.720 ;
        RECT 69.590 33.550 69.760 33.720 ;
        RECT 69.950 33.550 70.120 33.720 ;
        RECT 21.905 32.620 22.075 32.790 ;
        RECT 22.265 32.620 22.435 32.790 ;
        RECT 22.625 32.620 22.795 32.790 ;
        RECT 22.985 32.620 23.155 32.790 ;
        RECT 23.345 32.620 23.515 32.790 ;
        RECT 23.705 32.620 23.875 32.790 ;
        RECT 34.900 32.620 35.070 32.790 ;
        RECT 35.260 32.620 35.430 32.790 ;
        RECT 35.620 32.620 35.790 32.790 ;
        RECT 35.980 32.620 36.150 32.790 ;
        RECT 36.340 32.620 36.510 32.790 ;
        RECT 36.700 32.620 36.870 32.790 ;
        RECT 40.325 32.405 40.495 32.575 ;
        RECT 41.385 32.405 41.555 32.575 ;
        RECT 43.715 32.405 43.885 32.575 ;
        RECT 48.570 32.690 48.740 32.860 ;
        RECT 51.570 32.690 51.740 32.860 ;
        RECT 55.155 32.720 55.325 32.890 ;
        RECT 55.515 32.720 55.685 32.890 ;
        RECT 55.875 32.720 56.045 32.890 ;
        RECT 56.235 32.720 56.405 32.890 ;
        RECT 56.595 32.720 56.765 32.890 ;
        RECT 56.955 32.720 57.125 32.890 ;
        RECT 68.150 32.720 68.320 32.890 ;
        RECT 68.510 32.720 68.680 32.890 ;
        RECT 68.870 32.720 69.040 32.890 ;
        RECT 69.230 32.720 69.400 32.890 ;
        RECT 69.590 32.720 69.760 32.890 ;
        RECT 69.950 32.720 70.120 32.890 ;
        RECT 44.775 32.405 44.945 32.575 ;
        RECT 48.085 32.295 48.255 32.465 ;
        RECT 21.905 31.790 22.075 31.960 ;
        RECT 22.265 31.790 22.435 31.960 ;
        RECT 22.625 31.790 22.795 31.960 ;
        RECT 22.985 31.790 23.155 31.960 ;
        RECT 23.345 31.790 23.515 31.960 ;
        RECT 23.705 31.790 23.875 31.960 ;
        RECT 40.855 32.010 41.025 32.180 ;
        RECT 44.245 32.010 44.415 32.180 ;
        RECT 49.055 32.295 49.225 32.465 ;
        RECT 51.085 32.295 51.255 32.465 ;
        RECT 52.055 32.295 52.225 32.465 ;
        RECT 34.900 31.790 35.070 31.960 ;
        RECT 35.260 31.790 35.430 31.960 ;
        RECT 35.620 31.790 35.790 31.960 ;
        RECT 35.980 31.790 36.150 31.960 ;
        RECT 36.340 31.790 36.510 31.960 ;
        RECT 36.700 31.790 36.870 31.960 ;
        RECT 48.570 31.900 48.740 32.070 ;
        RECT 55.155 31.890 55.325 32.060 ;
        RECT 55.515 31.890 55.685 32.060 ;
        RECT 55.875 31.890 56.045 32.060 ;
        RECT 56.235 31.890 56.405 32.060 ;
        RECT 56.595 31.890 56.765 32.060 ;
        RECT 56.955 31.890 57.125 32.060 ;
        RECT 68.150 31.890 68.320 32.060 ;
        RECT 68.510 31.890 68.680 32.060 ;
        RECT 68.870 31.890 69.040 32.060 ;
        RECT 69.230 31.890 69.400 32.060 ;
        RECT 69.590 31.890 69.760 32.060 ;
        RECT 69.950 31.890 70.120 32.060 ;
        RECT 21.905 30.960 22.075 31.130 ;
        RECT 22.265 30.960 22.435 31.130 ;
        RECT 22.625 30.960 22.795 31.130 ;
        RECT 22.985 30.960 23.155 31.130 ;
        RECT 23.345 30.960 23.515 31.130 ;
        RECT 23.705 30.960 23.875 31.130 ;
        RECT 34.900 30.960 35.070 31.130 ;
        RECT 35.260 30.960 35.430 31.130 ;
        RECT 35.620 30.960 35.790 31.130 ;
        RECT 35.980 30.960 36.150 31.130 ;
        RECT 36.340 30.960 36.510 31.130 ;
        RECT 36.700 30.960 36.870 31.130 ;
        RECT 55.155 31.060 55.325 31.230 ;
        RECT 55.515 31.060 55.685 31.230 ;
        RECT 55.875 31.060 56.045 31.230 ;
        RECT 56.235 31.060 56.405 31.230 ;
        RECT 56.595 31.060 56.765 31.230 ;
        RECT 56.955 31.060 57.125 31.230 ;
        RECT 68.150 31.060 68.320 31.230 ;
        RECT 68.510 31.060 68.680 31.230 ;
        RECT 68.870 31.060 69.040 31.230 ;
        RECT 69.230 31.060 69.400 31.230 ;
        RECT 69.590 31.060 69.760 31.230 ;
        RECT 69.950 31.060 70.120 31.230 ;
        RECT 21.905 30.130 22.075 30.300 ;
        RECT 22.265 30.130 22.435 30.300 ;
        RECT 22.625 30.130 22.795 30.300 ;
        RECT 22.985 30.130 23.155 30.300 ;
        RECT 23.345 30.130 23.515 30.300 ;
        RECT 23.705 30.130 23.875 30.300 ;
        RECT 34.900 30.130 35.070 30.300 ;
        RECT 35.260 30.130 35.430 30.300 ;
        RECT 35.620 30.130 35.790 30.300 ;
        RECT 35.980 30.130 36.150 30.300 ;
        RECT 36.340 30.130 36.510 30.300 ;
        RECT 36.700 30.130 36.870 30.300 ;
        RECT 55.155 30.230 55.325 30.400 ;
        RECT 55.515 30.230 55.685 30.400 ;
        RECT 55.875 30.230 56.045 30.400 ;
        RECT 56.235 30.230 56.405 30.400 ;
        RECT 56.595 30.230 56.765 30.400 ;
        RECT 56.955 30.230 57.125 30.400 ;
        RECT 68.150 30.230 68.320 30.400 ;
        RECT 68.510 30.230 68.680 30.400 ;
        RECT 68.870 30.230 69.040 30.400 ;
        RECT 69.230 30.230 69.400 30.400 ;
        RECT 69.590 30.230 69.760 30.400 ;
        RECT 69.950 30.230 70.120 30.400 ;
        RECT 48.580 29.910 48.750 30.080 ;
        RECT 51.570 29.910 51.740 30.080 ;
        RECT 21.905 29.300 22.075 29.470 ;
        RECT 22.265 29.300 22.435 29.470 ;
        RECT 22.625 29.300 22.795 29.470 ;
        RECT 22.985 29.300 23.155 29.470 ;
        RECT 23.345 29.300 23.515 29.470 ;
        RECT 23.705 29.300 23.875 29.470 ;
        RECT 34.900 29.300 35.070 29.470 ;
        RECT 35.260 29.300 35.430 29.470 ;
        RECT 35.620 29.300 35.790 29.470 ;
        RECT 35.980 29.300 36.150 29.470 ;
        RECT 36.340 29.300 36.510 29.470 ;
        RECT 36.700 29.300 36.870 29.470 ;
        RECT 48.095 29.515 48.265 29.685 ;
        RECT 49.065 29.515 49.235 29.685 ;
        RECT 51.085 29.515 51.255 29.685 ;
        RECT 52.055 29.515 52.225 29.685 ;
        RECT 55.155 29.400 55.325 29.570 ;
        RECT 55.515 29.400 55.685 29.570 ;
        RECT 55.875 29.400 56.045 29.570 ;
        RECT 56.235 29.400 56.405 29.570 ;
        RECT 56.595 29.400 56.765 29.570 ;
        RECT 56.955 29.400 57.125 29.570 ;
        RECT 68.150 29.400 68.320 29.570 ;
        RECT 68.510 29.400 68.680 29.570 ;
        RECT 68.870 29.400 69.040 29.570 ;
        RECT 69.230 29.400 69.400 29.570 ;
        RECT 69.590 29.400 69.760 29.570 ;
        RECT 69.950 29.400 70.120 29.570 ;
        RECT 48.580 29.120 48.750 29.290 ;
        RECT 21.905 28.470 22.075 28.640 ;
        RECT 22.265 28.470 22.435 28.640 ;
        RECT 22.625 28.470 22.795 28.640 ;
        RECT 22.985 28.470 23.155 28.640 ;
        RECT 23.345 28.470 23.515 28.640 ;
        RECT 23.705 28.470 23.875 28.640 ;
        RECT 34.900 28.470 35.070 28.640 ;
        RECT 35.260 28.470 35.430 28.640 ;
        RECT 35.620 28.470 35.790 28.640 ;
        RECT 35.980 28.470 36.150 28.640 ;
        RECT 36.340 28.470 36.510 28.640 ;
        RECT 36.700 28.470 36.870 28.640 ;
        RECT 55.155 28.570 55.325 28.740 ;
        RECT 55.515 28.570 55.685 28.740 ;
        RECT 55.875 28.570 56.045 28.740 ;
        RECT 56.235 28.570 56.405 28.740 ;
        RECT 56.595 28.570 56.765 28.740 ;
        RECT 56.955 28.570 57.125 28.740 ;
        RECT 68.150 28.570 68.320 28.740 ;
        RECT 68.510 28.570 68.680 28.740 ;
        RECT 68.870 28.570 69.040 28.740 ;
        RECT 69.230 28.570 69.400 28.740 ;
        RECT 69.590 28.570 69.760 28.740 ;
        RECT 69.950 28.570 70.120 28.740 ;
        RECT 21.905 27.640 22.075 27.810 ;
        RECT 22.265 27.640 22.435 27.810 ;
        RECT 22.625 27.640 22.795 27.810 ;
        RECT 22.985 27.640 23.155 27.810 ;
        RECT 23.345 27.640 23.515 27.810 ;
        RECT 23.705 27.640 23.875 27.810 ;
        RECT 34.900 27.640 35.070 27.810 ;
        RECT 35.260 27.640 35.430 27.810 ;
        RECT 35.620 27.640 35.790 27.810 ;
        RECT 35.980 27.640 36.150 27.810 ;
        RECT 36.340 27.640 36.510 27.810 ;
        RECT 36.700 27.640 36.870 27.810 ;
        RECT 55.155 27.740 55.325 27.910 ;
        RECT 55.515 27.740 55.685 27.910 ;
        RECT 55.875 27.740 56.045 27.910 ;
        RECT 56.235 27.740 56.405 27.910 ;
        RECT 56.595 27.740 56.765 27.910 ;
        RECT 56.955 27.740 57.125 27.910 ;
        RECT 68.150 27.740 68.320 27.910 ;
        RECT 68.510 27.740 68.680 27.910 ;
        RECT 68.870 27.740 69.040 27.910 ;
        RECT 69.230 27.740 69.400 27.910 ;
        RECT 69.590 27.740 69.760 27.910 ;
        RECT 69.950 27.740 70.120 27.910 ;
        RECT 48.580 27.130 48.750 27.300 ;
        RECT 21.905 26.810 22.075 26.980 ;
        RECT 22.265 26.810 22.435 26.980 ;
        RECT 22.625 26.810 22.795 26.980 ;
        RECT 22.985 26.810 23.155 26.980 ;
        RECT 23.345 26.810 23.515 26.980 ;
        RECT 23.705 26.810 23.875 26.980 ;
        RECT 34.900 26.810 35.070 26.980 ;
        RECT 35.260 26.810 35.430 26.980 ;
        RECT 35.620 26.810 35.790 26.980 ;
        RECT 35.980 26.810 36.150 26.980 ;
        RECT 36.340 26.810 36.510 26.980 ;
        RECT 36.700 26.810 36.870 26.980 ;
        RECT 48.095 26.735 48.265 26.905 ;
        RECT 49.065 26.735 49.235 26.905 ;
        RECT 55.155 26.910 55.325 27.080 ;
        RECT 55.515 26.910 55.685 27.080 ;
        RECT 55.875 26.910 56.045 27.080 ;
        RECT 56.235 26.910 56.405 27.080 ;
        RECT 56.595 26.910 56.765 27.080 ;
        RECT 56.955 26.910 57.125 27.080 ;
        RECT 68.150 26.910 68.320 27.080 ;
        RECT 68.510 26.910 68.680 27.080 ;
        RECT 68.870 26.910 69.040 27.080 ;
        RECT 69.230 26.910 69.400 27.080 ;
        RECT 69.590 26.910 69.760 27.080 ;
        RECT 69.950 26.910 70.120 27.080 ;
        RECT 21.905 25.980 22.075 26.150 ;
        RECT 22.265 25.980 22.435 26.150 ;
        RECT 22.625 25.980 22.795 26.150 ;
        RECT 22.985 25.980 23.155 26.150 ;
        RECT 23.345 25.980 23.515 26.150 ;
        RECT 23.705 25.980 23.875 26.150 ;
        RECT 34.900 25.980 35.070 26.150 ;
        RECT 35.260 25.980 35.430 26.150 ;
        RECT 35.620 25.980 35.790 26.150 ;
        RECT 35.980 25.980 36.150 26.150 ;
        RECT 36.340 25.980 36.510 26.150 ;
        RECT 36.700 25.980 36.870 26.150 ;
        RECT 55.155 26.080 55.325 26.250 ;
        RECT 55.515 26.080 55.685 26.250 ;
        RECT 55.875 26.080 56.045 26.250 ;
        RECT 56.235 26.080 56.405 26.250 ;
        RECT 56.595 26.080 56.765 26.250 ;
        RECT 56.955 26.080 57.125 26.250 ;
        RECT 68.150 26.080 68.320 26.250 ;
        RECT 68.510 26.080 68.680 26.250 ;
        RECT 68.870 26.080 69.040 26.250 ;
        RECT 69.230 26.080 69.400 26.250 ;
        RECT 69.590 26.080 69.760 26.250 ;
        RECT 69.950 26.080 70.120 26.250 ;
        RECT 21.905 25.150 22.075 25.320 ;
        RECT 22.265 25.150 22.435 25.320 ;
        RECT 22.625 25.150 22.795 25.320 ;
        RECT 22.985 25.150 23.155 25.320 ;
        RECT 23.345 25.150 23.515 25.320 ;
        RECT 23.705 25.150 23.875 25.320 ;
        RECT 34.900 25.150 35.070 25.320 ;
        RECT 35.260 25.150 35.430 25.320 ;
        RECT 35.620 25.150 35.790 25.320 ;
        RECT 35.980 25.150 36.150 25.320 ;
        RECT 36.340 25.150 36.510 25.320 ;
        RECT 36.700 25.150 36.870 25.320 ;
        RECT 55.155 25.250 55.325 25.420 ;
        RECT 55.515 25.250 55.685 25.420 ;
        RECT 55.875 25.250 56.045 25.420 ;
        RECT 56.235 25.250 56.405 25.420 ;
        RECT 56.595 25.250 56.765 25.420 ;
        RECT 56.955 25.250 57.125 25.420 ;
        RECT 68.150 25.250 68.320 25.420 ;
        RECT 68.510 25.250 68.680 25.420 ;
        RECT 68.870 25.250 69.040 25.420 ;
        RECT 69.230 25.250 69.400 25.420 ;
        RECT 69.590 25.250 69.760 25.420 ;
        RECT 69.950 25.250 70.120 25.420 ;
        RECT 21.905 24.320 22.075 24.490 ;
        RECT 22.265 24.320 22.435 24.490 ;
        RECT 22.625 24.320 22.795 24.490 ;
        RECT 22.985 24.320 23.155 24.490 ;
        RECT 23.345 24.320 23.515 24.490 ;
        RECT 23.705 24.320 23.875 24.490 ;
        RECT 34.900 24.320 35.070 24.490 ;
        RECT 35.260 24.320 35.430 24.490 ;
        RECT 35.620 24.320 35.790 24.490 ;
        RECT 35.980 24.320 36.150 24.490 ;
        RECT 36.340 24.320 36.510 24.490 ;
        RECT 36.700 24.320 36.870 24.490 ;
        RECT 55.155 24.420 55.325 24.590 ;
        RECT 55.515 24.420 55.685 24.590 ;
        RECT 55.875 24.420 56.045 24.590 ;
        RECT 56.235 24.420 56.405 24.590 ;
        RECT 56.595 24.420 56.765 24.590 ;
        RECT 56.955 24.420 57.125 24.590 ;
        RECT 68.150 24.420 68.320 24.590 ;
        RECT 68.510 24.420 68.680 24.590 ;
        RECT 68.870 24.420 69.040 24.590 ;
        RECT 69.230 24.420 69.400 24.590 ;
        RECT 69.590 24.420 69.760 24.590 ;
        RECT 69.950 24.420 70.120 24.590 ;
        RECT 21.905 23.490 22.075 23.660 ;
        RECT 22.265 23.490 22.435 23.660 ;
        RECT 22.625 23.490 22.795 23.660 ;
        RECT 22.985 23.490 23.155 23.660 ;
        RECT 23.345 23.490 23.515 23.660 ;
        RECT 23.705 23.490 23.875 23.660 ;
        RECT 34.900 23.490 35.070 23.660 ;
        RECT 35.260 23.490 35.430 23.660 ;
        RECT 35.620 23.490 35.790 23.660 ;
        RECT 35.980 23.490 36.150 23.660 ;
        RECT 36.340 23.490 36.510 23.660 ;
        RECT 36.700 23.490 36.870 23.660 ;
        RECT 55.155 23.590 55.325 23.760 ;
        RECT 55.515 23.590 55.685 23.760 ;
        RECT 55.875 23.590 56.045 23.760 ;
        RECT 56.235 23.590 56.405 23.760 ;
        RECT 56.595 23.590 56.765 23.760 ;
        RECT 56.955 23.590 57.125 23.760 ;
        RECT 68.150 23.590 68.320 23.760 ;
        RECT 68.510 23.590 68.680 23.760 ;
        RECT 68.870 23.590 69.040 23.760 ;
        RECT 69.230 23.590 69.400 23.760 ;
        RECT 69.590 23.590 69.760 23.760 ;
        RECT 69.950 23.590 70.120 23.760 ;
        RECT 21.905 22.660 22.075 22.830 ;
        RECT 22.265 22.660 22.435 22.830 ;
        RECT 22.625 22.660 22.795 22.830 ;
        RECT 22.985 22.660 23.155 22.830 ;
        RECT 23.345 22.660 23.515 22.830 ;
        RECT 23.705 22.660 23.875 22.830 ;
        RECT 34.900 22.660 35.070 22.830 ;
        RECT 35.260 22.660 35.430 22.830 ;
        RECT 35.620 22.660 35.790 22.830 ;
        RECT 35.980 22.660 36.150 22.830 ;
        RECT 36.340 22.660 36.510 22.830 ;
        RECT 36.700 22.660 36.870 22.830 ;
        RECT 68.150 22.760 68.320 22.930 ;
        RECT 68.510 22.760 68.680 22.930 ;
        RECT 68.870 22.760 69.040 22.930 ;
        RECT 69.230 22.760 69.400 22.930 ;
        RECT 69.590 22.760 69.760 22.930 ;
        RECT 69.950 22.760 70.120 22.930 ;
      LAYER met1 ;
        RECT 43.115 80.060 47.855 80.300 ;
        RECT 43.115 79.930 43.355 80.060 ;
        RECT 42.585 79.690 43.355 79.930 ;
        RECT 47.615 79.935 47.855 80.060 ;
        RECT 47.615 79.745 48.875 79.935 ;
        RECT 47.615 79.695 48.930 79.745 ;
        RECT 42.610 79.480 43.110 79.690 ;
        RECT 43.270 79.295 43.660 79.520 ;
        RECT 45.425 79.295 45.655 79.535 ;
        RECT 48.430 79.515 48.930 79.695 ;
        RECT 43.270 79.245 45.655 79.295 ;
        RECT 43.270 79.230 45.650 79.245 ;
        RECT 43.390 79.090 45.650 79.230 ;
        RECT 21.805 77.350 23.965 78.530 ;
        RECT 34.770 78.290 39.670 78.665 ;
        RECT 44.490 78.425 44.735 79.090 ;
        RECT 34.830 78.230 36.935 78.290 ;
        RECT 21.805 75.690 23.965 76.870 ;
        RECT 34.805 76.520 36.965 77.700 ;
        RECT 21.805 74.030 23.965 75.210 ;
        RECT 34.805 74.860 36.965 76.040 ;
        RECT 21.805 72.370 23.965 73.550 ;
        RECT 34.805 73.200 36.965 74.380 ;
        RECT 39.295 72.845 39.670 78.290 ;
        RECT 44.445 77.445 44.805 78.425 ;
        RECT 44.530 77.330 44.805 77.445 ;
        RECT 52.150 78.290 57.230 78.665 ;
        RECT 44.530 77.140 46.545 77.330 ;
        RECT 46.355 76.880 46.545 77.140 ;
        RECT 46.690 76.880 47.110 76.905 ;
        RECT 46.355 76.690 47.125 76.880 ;
        RECT 46.690 76.675 47.110 76.690 ;
        RECT 43.565 75.140 44.565 75.320 ;
        RECT 46.755 75.140 47.755 75.320 ;
        RECT 43.565 75.090 47.785 75.140 ;
        RECT 43.935 74.930 47.785 75.090 ;
        RECT 43.965 74.440 44.295 74.930 ;
        RECT 52.150 72.845 52.525 78.290 ;
        RECT 55.055 76.620 57.215 77.800 ;
        RECT 68.055 77.450 70.215 78.630 ;
        RECT 55.055 74.960 57.215 76.140 ;
        RECT 68.055 75.790 70.215 76.970 ;
        RECT 55.055 73.300 57.215 74.480 ;
        RECT 68.055 74.130 70.215 75.310 ;
        RECT 21.805 70.710 23.965 71.890 ;
        RECT 34.805 71.540 36.965 72.720 ;
        RECT 39.295 72.470 52.525 72.845 ;
        RECT 42.455 71.920 42.685 71.980 ;
        RECT 43.905 71.920 44.265 72.180 ;
        RECT 42.455 71.760 44.265 71.920 ;
        RECT 42.455 71.690 42.685 71.760 ;
        RECT 43.905 71.200 44.265 71.760 ;
        RECT 55.055 71.640 57.215 72.820 ;
        RECT 68.055 72.470 70.215 73.650 ;
        RECT 21.805 69.050 23.965 70.230 ;
        RECT 34.805 69.880 36.965 71.060 ;
        RECT 55.055 69.980 57.215 71.160 ;
        RECT 68.055 70.810 70.215 71.990 ;
        RECT 21.805 67.390 23.965 68.570 ;
        RECT 34.805 68.220 36.965 69.400 ;
        RECT 55.055 68.320 57.215 69.500 ;
        RECT 68.055 69.150 70.215 70.330 ;
        RECT 21.805 65.730 23.965 66.910 ;
        RECT 34.805 66.560 36.965 67.740 ;
        RECT 45.745 67.700 49.505 67.980 ;
        RECT 45.745 67.650 49.510 67.700 ;
        RECT 45.750 67.440 46.170 67.650 ;
        RECT 49.090 67.470 49.510 67.650 ;
        RECT 45.315 67.250 45.545 67.390 ;
        RECT 46.355 67.250 46.685 67.450 ;
        RECT 48.655 67.320 48.885 67.420 ;
        RECT 49.715 67.320 49.945 67.420 ;
        RECT 45.315 67.040 46.685 67.250 ;
        RECT 45.315 66.930 45.545 67.040 ;
        RECT 42.235 66.700 42.655 66.870 ;
        RECT 45.255 66.700 45.585 66.750 ;
        RECT 45.750 66.700 46.170 66.880 ;
        RECT 46.355 66.860 46.685 67.040 ;
        RECT 48.165 67.060 49.945 67.320 ;
        RECT 47.005 66.700 47.335 66.760 ;
        RECT 48.165 66.700 48.425 67.060 ;
        RECT 48.655 66.960 48.885 67.060 ;
        RECT 49.715 66.960 49.945 67.060 ;
        RECT 42.225 66.440 48.425 66.700 ;
        RECT 55.055 66.660 57.215 67.840 ;
        RECT 68.055 67.490 70.215 68.670 ;
        RECT 45.255 66.160 45.585 66.440 ;
        RECT 47.005 66.170 47.335 66.440 ;
        RECT 21.805 64.070 23.965 65.250 ;
        RECT 34.805 64.900 36.965 66.080 ;
        RECT 46.345 64.850 46.675 65.110 ;
        RECT 48.125 64.850 48.455 65.110 ;
        RECT 55.055 65.000 57.215 66.180 ;
        RECT 68.055 65.830 70.215 67.010 ;
        RECT 42.205 64.590 48.455 64.850 ;
        RECT 21.805 62.410 23.965 63.590 ;
        RECT 34.805 63.240 36.965 64.420 ;
        RECT 42.245 64.400 42.665 64.590 ;
        RECT 41.855 64.220 42.085 64.350 ;
        RECT 42.825 64.220 43.055 64.350 ;
        RECT 43.965 64.220 44.295 64.390 ;
        RECT 41.855 64.020 44.295 64.220 ;
        RECT 41.855 63.890 42.085 64.020 ;
        RECT 42.825 63.890 43.055 64.020 ;
        RECT 43.965 63.800 44.295 64.020 ;
        RECT 45.255 64.250 45.585 64.400 ;
        RECT 45.740 64.390 46.160 64.590 ;
        RECT 46.345 64.520 46.675 64.590 ;
        RECT 48.125 64.520 48.455 64.590 ;
        RECT 46.365 64.250 46.595 64.340 ;
        RECT 45.255 64.040 46.675 64.250 ;
        RECT 48.155 64.230 48.415 64.520 ;
        RECT 48.655 64.230 48.885 64.340 ;
        RECT 49.715 64.230 49.945 64.340 ;
        RECT 45.255 63.810 45.585 64.040 ;
        RECT 46.365 63.880 46.595 64.040 ;
        RECT 48.155 63.970 49.945 64.230 ;
        RECT 48.655 63.880 48.885 63.970 ;
        RECT 49.715 63.880 49.945 63.970 ;
        RECT 21.805 60.750 23.965 61.930 ;
        RECT 34.805 61.580 36.965 62.760 ;
        RECT 44.005 62.380 44.245 63.800 ;
        RECT 45.740 63.640 46.160 63.830 ;
        RECT 49.090 63.640 49.510 63.830 ;
        RECT 45.740 63.600 49.510 63.640 ;
        RECT 45.745 63.310 49.505 63.600 ;
        RECT 55.055 63.340 57.215 64.520 ;
        RECT 68.055 64.170 70.215 65.350 ;
        RECT 47.015 62.380 47.345 63.110 ;
        RECT 48.165 62.410 48.495 63.110 ;
        RECT 43.695 61.380 44.695 62.380 ;
        RECT 46.385 61.380 47.385 62.380 ;
        RECT 48.125 61.410 49.125 62.410 ;
        RECT 55.055 61.680 57.215 62.860 ;
        RECT 68.055 62.510 70.215 63.690 ;
        RECT 21.805 59.090 23.965 60.270 ;
        RECT 34.805 59.920 36.965 61.100 ;
        RECT 42.865 60.100 43.255 61.155 ;
        RECT 46.910 60.420 47.080 61.380 ;
        RECT 48.000 60.420 48.320 60.685 ;
        RECT 46.910 60.250 48.320 60.420 ;
        RECT 21.805 57.430 23.965 58.610 ;
        RECT 34.805 58.260 36.965 59.440 ;
        RECT 42.970 58.980 43.160 60.100 ;
        RECT 48.000 59.650 48.320 60.250 ;
        RECT 55.055 60.020 57.215 61.200 ;
        RECT 68.055 60.850 70.215 62.030 ;
        RECT 42.970 58.790 48.880 58.980 ;
        RECT 49.690 58.850 51.855 58.975 ;
        RECT 44.120 58.680 44.540 58.790 ;
        RECT 43.685 58.500 43.915 58.630 ;
        RECT 44.745 58.500 44.975 58.630 ;
        RECT 48.455 58.620 48.875 58.790 ;
        RECT 49.690 58.785 51.875 58.850 ;
        RECT 43.685 58.280 45.460 58.500 ;
        RECT 43.685 58.170 43.915 58.280 ;
        RECT 44.745 58.170 44.975 58.280 ;
        RECT 21.805 55.770 23.965 56.950 ;
        RECT 34.805 56.600 36.965 57.780 ;
        RECT 45.240 56.235 45.460 58.280 ;
        RECT 48.455 57.910 48.875 58.060 ;
        RECT 49.690 57.910 49.880 58.785 ;
        RECT 51.455 58.620 51.875 58.785 ;
        RECT 51.065 58.450 51.295 58.570 ;
        RECT 52.035 58.450 52.265 58.570 ;
        RECT 48.455 57.830 49.880 57.910 ;
        RECT 48.505 57.720 49.880 57.830 ;
        RECT 50.570 58.230 52.265 58.450 ;
        RECT 55.055 58.360 57.215 59.540 ;
        RECT 68.055 59.190 70.215 60.370 ;
        RECT 50.570 56.305 50.790 58.230 ;
        RECT 51.065 58.110 51.295 58.230 ;
        RECT 52.035 58.110 52.265 58.230 ;
        RECT 55.055 56.700 57.215 57.880 ;
        RECT 68.055 57.530 70.215 58.710 ;
        RECT 50.570 56.235 50.785 56.305 ;
        RECT 21.805 54.110 23.965 55.290 ;
        RECT 34.805 54.940 36.965 56.120 ;
        RECT 45.240 56.015 50.785 56.235 ;
        RECT 46.355 54.845 46.690 56.015 ;
        RECT 55.055 55.040 57.215 56.220 ;
        RECT 68.055 55.870 70.215 57.050 ;
        RECT 46.145 54.720 46.970 54.845 ;
        RECT 44.085 54.525 47.840 54.720 ;
        RECT 21.805 52.450 23.965 53.630 ;
        RECT 34.805 53.280 36.965 54.460 ;
        RECT 44.120 54.330 44.540 54.525 ;
        RECT 46.145 54.460 46.970 54.525 ;
        RECT 40.195 54.280 40.430 54.310 ;
        RECT 40.195 54.130 40.525 54.280 ;
        RECT 41.355 54.130 41.585 54.280 ;
        RECT 40.195 53.975 41.585 54.130 ;
        RECT 40.195 53.820 40.525 53.975 ;
        RECT 41.355 53.820 41.585 53.975 ;
        RECT 43.685 54.135 43.915 54.280 ;
        RECT 44.745 54.135 44.975 54.280 ;
        RECT 43.685 53.940 46.360 54.135 ;
        RECT 43.685 53.820 43.915 53.940 ;
        RECT 44.745 53.820 44.975 53.940 ;
        RECT 21.805 50.790 23.965 51.970 ;
        RECT 34.805 51.620 36.965 52.800 ;
        RECT 40.195 51.200 40.430 53.820 ;
        RECT 40.730 53.625 41.150 53.770 ;
        RECT 44.120 53.625 44.540 53.770 ;
        RECT 40.695 53.405 44.540 53.625 ;
        RECT 46.165 51.955 46.360 53.940 ;
        RECT 47.645 52.480 47.840 54.525 ;
        RECT 55.055 53.380 57.215 54.560 ;
        RECT 68.055 54.210 70.215 55.390 ;
        RECT 47.645 52.285 48.870 52.480 ;
        RECT 48.445 52.120 48.865 52.285 ;
        RECT 49.400 52.265 51.865 52.475 ;
        RECT 48.055 51.955 48.285 52.070 ;
        RECT 49.025 51.955 49.255 52.070 ;
        RECT 46.165 51.760 49.255 51.955 ;
        RECT 46.165 51.610 46.360 51.760 ;
        RECT 48.055 51.610 48.285 51.760 ;
        RECT 49.025 51.610 49.255 51.760 ;
        RECT 44.100 51.415 47.865 51.610 ;
        RECT 44.120 51.250 44.540 51.415 ;
        RECT 21.805 49.130 23.965 50.310 ;
        RECT 34.805 49.960 36.965 51.140 ;
        RECT 40.195 51.050 40.525 51.200 ;
        RECT 41.355 51.050 41.585 51.200 ;
        RECT 40.195 50.895 41.585 51.050 ;
        RECT 40.195 50.740 40.525 50.895 ;
        RECT 41.355 50.740 41.585 50.895 ;
        RECT 43.685 51.055 43.915 51.200 ;
        RECT 44.745 51.055 44.975 51.200 ;
        RECT 43.685 50.860 46.360 51.055 ;
        RECT 43.685 50.740 43.915 50.860 ;
        RECT 44.745 50.740 44.975 50.860 ;
        RECT 21.805 47.470 23.965 48.650 ;
        RECT 34.805 48.300 36.965 49.480 ;
        RECT 40.195 48.120 40.430 50.740 ;
        RECT 40.730 50.545 41.150 50.690 ;
        RECT 44.120 50.545 44.540 50.690 ;
        RECT 40.695 50.325 44.540 50.545 ;
        RECT 45.225 49.370 45.675 50.520 ;
        RECT 45.315 48.555 45.595 49.370 ;
        RECT 46.165 49.175 46.360 50.860 ;
        RECT 47.670 49.745 47.865 51.415 ;
        RECT 48.445 51.410 48.865 51.560 ;
        RECT 49.400 51.410 49.610 52.265 ;
        RECT 51.445 52.120 51.865 52.265 ;
        RECT 51.055 51.930 51.285 52.070 ;
        RECT 52.025 52.020 52.255 52.070 ;
        RECT 52.025 51.930 52.400 52.020 ;
        RECT 51.055 51.765 52.400 51.930 ;
        RECT 51.055 51.610 51.285 51.765 ;
        RECT 52.025 51.610 52.400 51.765 ;
        RECT 55.055 51.720 57.215 52.900 ;
        RECT 68.055 52.550 70.215 53.730 ;
        RECT 48.435 51.200 49.610 51.410 ;
        RECT 47.670 49.550 48.875 49.745 ;
        RECT 48.445 49.340 48.865 49.550 ;
        RECT 49.400 49.485 51.865 49.695 ;
        RECT 48.055 49.175 48.285 49.290 ;
        RECT 49.025 49.175 49.255 49.290 ;
        RECT 46.165 48.980 49.255 49.175 ;
        RECT 46.165 48.555 46.360 48.980 ;
        RECT 48.055 48.830 48.285 48.980 ;
        RECT 49.025 48.830 49.255 48.980 ;
        RECT 48.445 48.630 48.865 48.780 ;
        RECT 49.400 48.630 49.610 49.485 ;
        RECT 51.445 49.340 51.865 49.485 ;
        RECT 52.160 49.290 52.400 51.610 ;
        RECT 55.055 50.060 57.215 51.240 ;
        RECT 68.055 50.890 70.215 52.070 ;
        RECT 51.055 49.150 51.285 49.290 ;
        RECT 52.025 49.150 52.400 49.290 ;
        RECT 51.055 48.985 52.400 49.150 ;
        RECT 51.055 48.830 51.285 48.985 ;
        RECT 52.025 48.830 52.400 48.985 ;
        RECT 44.085 48.360 47.900 48.555 ;
        RECT 48.435 48.420 49.610 48.630 ;
        RECT 44.120 48.170 44.540 48.360 ;
        RECT 40.195 47.970 40.525 48.120 ;
        RECT 41.355 47.970 41.585 48.120 ;
        RECT 21.805 45.810 23.965 46.990 ;
        RECT 34.805 46.640 36.965 47.820 ;
        RECT 40.195 47.815 41.585 47.970 ;
        RECT 40.195 47.660 40.525 47.815 ;
        RECT 41.355 47.660 41.585 47.815 ;
        RECT 43.685 47.975 43.915 48.120 ;
        RECT 44.745 47.975 44.975 48.120 ;
        RECT 43.685 47.780 46.360 47.975 ;
        RECT 43.685 47.660 43.915 47.780 ;
        RECT 44.745 47.660 44.975 47.780 ;
        RECT 21.805 44.150 23.965 45.330 ;
        RECT 34.805 44.980 36.965 46.160 ;
        RECT 40.195 45.040 40.430 47.660 ;
        RECT 40.730 47.465 41.150 47.610 ;
        RECT 44.120 47.465 44.540 47.610 ;
        RECT 40.695 47.245 44.540 47.465 ;
        RECT 45.225 45.435 45.675 46.455 ;
        RECT 46.165 46.395 46.360 47.780 ;
        RECT 47.705 46.930 47.900 48.360 ;
        RECT 47.705 46.735 48.895 46.930 ;
        RECT 48.445 46.560 48.865 46.735 ;
        RECT 49.400 46.705 51.865 46.915 ;
        RECT 48.055 46.395 48.285 46.510 ;
        RECT 49.025 46.395 49.255 46.510 ;
        RECT 46.165 46.200 49.255 46.395 ;
        RECT 46.165 45.435 46.360 46.200 ;
        RECT 48.055 46.050 48.285 46.200 ;
        RECT 49.025 46.050 49.255 46.200 ;
        RECT 48.445 45.850 48.865 46.000 ;
        RECT 49.400 45.850 49.610 46.705 ;
        RECT 51.445 46.560 51.865 46.705 ;
        RECT 52.160 46.510 52.400 48.830 ;
        RECT 55.055 48.400 57.215 49.580 ;
        RECT 68.055 49.230 70.215 50.410 ;
        RECT 55.055 46.740 57.215 47.920 ;
        RECT 68.055 47.570 70.215 48.750 ;
        RECT 51.055 46.370 51.285 46.510 ;
        RECT 52.025 46.370 52.400 46.510 ;
        RECT 51.055 46.205 52.400 46.370 ;
        RECT 51.055 46.050 51.285 46.205 ;
        RECT 52.025 46.050 52.400 46.205 ;
        RECT 48.435 45.640 49.610 45.850 ;
        RECT 44.120 45.240 47.895 45.435 ;
        RECT 44.120 45.090 44.540 45.240 ;
        RECT 40.195 44.890 40.525 45.040 ;
        RECT 41.355 44.890 41.585 45.040 ;
        RECT 40.195 44.735 41.585 44.890 ;
        RECT 40.195 44.580 40.525 44.735 ;
        RECT 41.355 44.580 41.585 44.735 ;
        RECT 43.685 44.895 43.915 45.040 ;
        RECT 44.745 44.895 44.975 45.040 ;
        RECT 43.685 44.700 46.360 44.895 ;
        RECT 43.685 44.580 43.915 44.700 ;
        RECT 44.745 44.580 44.975 44.700 ;
        RECT 21.805 42.490 23.965 43.670 ;
        RECT 34.805 43.320 36.965 44.500 ;
        RECT 21.805 40.830 23.965 42.010 ;
        RECT 34.805 41.660 36.965 42.840 ;
        RECT 40.195 41.960 40.430 44.580 ;
        RECT 40.730 44.385 41.150 44.530 ;
        RECT 44.120 44.385 44.540 44.530 ;
        RECT 40.695 44.165 44.540 44.385 ;
        RECT 46.165 43.615 46.360 44.700 ;
        RECT 47.700 44.140 47.895 45.240 ;
        RECT 47.700 43.945 48.900 44.140 ;
        RECT 48.445 43.780 48.865 43.945 ;
        RECT 49.400 43.925 51.865 44.135 ;
        RECT 48.055 43.615 48.285 43.730 ;
        RECT 49.025 43.615 49.255 43.730 ;
        RECT 45.225 42.420 45.675 43.435 ;
        RECT 46.165 43.420 49.255 43.615 ;
        RECT 46.165 42.420 46.360 43.420 ;
        RECT 48.055 43.270 48.285 43.420 ;
        RECT 49.025 43.270 49.255 43.420 ;
        RECT 48.445 43.070 48.865 43.220 ;
        RECT 49.400 43.070 49.610 43.925 ;
        RECT 51.445 43.780 51.865 43.925 ;
        RECT 52.160 43.730 52.400 46.050 ;
        RECT 55.055 45.080 57.215 46.260 ;
        RECT 68.055 45.910 70.215 47.090 ;
        RECT 51.055 43.590 51.285 43.730 ;
        RECT 52.025 43.590 52.400 43.730 ;
        RECT 51.055 43.425 52.400 43.590 ;
        RECT 51.055 43.270 51.285 43.425 ;
        RECT 52.025 43.270 52.400 43.425 ;
        RECT 55.055 43.420 57.215 44.600 ;
        RECT 68.055 44.250 70.215 45.430 ;
        RECT 48.435 42.860 49.610 43.070 ;
        RECT 44.080 42.225 47.910 42.420 ;
        RECT 44.120 42.010 44.540 42.225 ;
        RECT 40.195 41.810 40.525 41.960 ;
        RECT 41.355 41.810 41.585 41.960 ;
        RECT 40.195 41.655 41.585 41.810 ;
        RECT 40.195 41.500 40.525 41.655 ;
        RECT 41.355 41.500 41.585 41.655 ;
        RECT 43.685 41.815 43.915 41.960 ;
        RECT 44.745 41.815 44.975 41.960 ;
        RECT 43.685 41.620 46.360 41.815 ;
        RECT 43.685 41.500 43.915 41.620 ;
        RECT 44.745 41.500 44.975 41.620 ;
        RECT 21.805 39.170 23.965 40.350 ;
        RECT 34.805 40.000 36.965 41.180 ;
        RECT 21.805 37.510 23.965 38.690 ;
        RECT 34.805 38.340 36.965 39.520 ;
        RECT 40.195 38.880 40.430 41.500 ;
        RECT 40.730 41.305 41.150 41.450 ;
        RECT 44.120 41.305 44.540 41.450 ;
        RECT 40.695 41.085 44.540 41.305 ;
        RECT 46.165 40.835 46.360 41.620 ;
        RECT 47.715 41.370 47.910 42.225 ;
        RECT 47.715 41.230 48.860 41.370 ;
        RECT 47.715 41.175 48.865 41.230 ;
        RECT 48.445 41.000 48.865 41.175 ;
        RECT 49.400 41.145 51.865 41.355 ;
        RECT 48.055 40.835 48.285 40.950 ;
        RECT 49.025 40.835 49.255 40.950 ;
        RECT 46.165 40.640 49.255 40.835 ;
        RECT 45.225 39.290 45.675 40.275 ;
        RECT 46.165 39.290 46.360 40.640 ;
        RECT 48.055 40.490 48.285 40.640 ;
        RECT 49.025 40.490 49.255 40.640 ;
        RECT 48.445 40.290 48.865 40.440 ;
        RECT 49.400 40.290 49.610 41.145 ;
        RECT 51.445 41.000 51.865 41.145 ;
        RECT 52.160 40.950 52.400 43.270 ;
        RECT 55.055 41.760 57.215 42.940 ;
        RECT 68.055 42.590 70.215 43.770 ;
        RECT 51.055 40.810 51.285 40.950 ;
        RECT 52.025 40.810 52.400 40.950 ;
        RECT 51.055 40.645 52.400 40.810 ;
        RECT 51.055 40.490 51.285 40.645 ;
        RECT 52.025 40.490 52.400 40.645 ;
        RECT 48.435 40.080 49.610 40.290 ;
        RECT 44.115 39.095 47.920 39.290 ;
        RECT 44.120 38.930 44.540 39.095 ;
        RECT 40.195 38.730 40.525 38.880 ;
        RECT 41.355 38.730 41.585 38.880 ;
        RECT 40.195 38.575 41.585 38.730 ;
        RECT 40.195 38.420 40.525 38.575 ;
        RECT 41.355 38.420 41.585 38.575 ;
        RECT 43.685 38.735 43.915 38.880 ;
        RECT 44.745 38.735 44.975 38.880 ;
        RECT 43.685 38.540 46.370 38.735 ;
        RECT 43.685 38.420 43.915 38.540 ;
        RECT 44.745 38.420 44.975 38.540 ;
        RECT 21.805 35.850 23.965 37.030 ;
        RECT 34.805 36.680 36.965 37.860 ;
        RECT 21.805 34.190 23.965 35.370 ;
        RECT 34.805 35.020 36.965 36.200 ;
        RECT 40.195 35.800 40.430 38.420 ;
        RECT 40.730 38.225 41.150 38.370 ;
        RECT 44.120 38.225 44.540 38.370 ;
        RECT 40.695 38.005 44.540 38.225 ;
        RECT 46.175 38.055 46.370 38.540 ;
        RECT 47.725 38.590 47.920 39.095 ;
        RECT 47.725 38.395 48.900 38.590 ;
        RECT 48.445 38.220 48.865 38.395 ;
        RECT 49.400 38.365 51.865 38.575 ;
        RECT 48.055 38.055 48.285 38.170 ;
        RECT 49.025 38.055 49.255 38.170 ;
        RECT 46.175 37.860 49.255 38.055 ;
        RECT 45.225 36.145 45.675 37.120 ;
        RECT 46.175 36.145 46.370 37.860 ;
        RECT 48.055 37.710 48.285 37.860 ;
        RECT 49.025 37.710 49.255 37.860 ;
        RECT 48.445 37.510 48.865 37.660 ;
        RECT 49.400 37.510 49.610 38.365 ;
        RECT 51.445 38.220 51.865 38.365 ;
        RECT 52.160 38.170 52.400 40.490 ;
        RECT 55.055 40.100 57.215 41.280 ;
        RECT 68.055 40.930 70.215 42.110 ;
        RECT 55.055 38.440 57.215 39.620 ;
        RECT 68.055 39.270 70.215 40.450 ;
        RECT 51.055 38.030 51.285 38.170 ;
        RECT 52.025 38.030 52.400 38.170 ;
        RECT 51.055 37.865 52.400 38.030 ;
        RECT 51.055 37.710 51.285 37.865 ;
        RECT 52.025 37.710 52.400 37.865 ;
        RECT 48.435 37.300 49.610 37.510 ;
        RECT 44.135 36.080 47.925 36.145 ;
        RECT 44.120 35.950 47.925 36.080 ;
        RECT 44.120 35.850 44.540 35.950 ;
        RECT 47.730 35.835 47.925 35.950 ;
        RECT 40.195 35.650 40.525 35.800 ;
        RECT 41.355 35.650 41.585 35.800 ;
        RECT 40.195 35.495 41.585 35.650 ;
        RECT 40.195 35.340 40.525 35.495 ;
        RECT 41.355 35.340 41.585 35.495 ;
        RECT 43.685 35.655 43.915 35.800 ;
        RECT 44.745 35.655 44.975 35.800 ;
        RECT 43.685 35.460 46.375 35.655 ;
        RECT 47.730 35.640 48.870 35.835 ;
        RECT 43.685 35.340 43.915 35.460 ;
        RECT 44.745 35.340 44.975 35.460 ;
        RECT 46.165 35.350 46.375 35.460 ;
        RECT 48.445 35.440 48.865 35.640 ;
        RECT 49.400 35.585 51.865 35.795 ;
        RECT 21.805 32.530 23.965 33.710 ;
        RECT 34.805 33.360 36.965 34.540 ;
        RECT 21.805 30.870 23.965 32.050 ;
        RECT 34.805 31.700 36.965 32.880 ;
        RECT 40.195 32.720 40.430 35.340 ;
        RECT 40.730 35.145 41.150 35.290 ;
        RECT 44.120 35.145 44.540 35.290 ;
        RECT 40.695 34.925 44.540 35.145 ;
        RECT 46.165 35.275 46.990 35.350 ;
        RECT 48.055 35.275 48.285 35.390 ;
        RECT 49.025 35.275 49.255 35.390 ;
        RECT 46.165 35.080 49.255 35.275 ;
        RECT 46.165 34.965 46.990 35.080 ;
        RECT 48.055 34.930 48.285 35.080 ;
        RECT 49.025 34.930 49.255 35.080 ;
        RECT 48.445 34.730 48.865 34.880 ;
        RECT 49.400 34.730 49.610 35.585 ;
        RECT 51.445 35.440 51.865 35.585 ;
        RECT 52.160 35.390 52.400 37.710 ;
        RECT 55.055 36.780 57.215 37.960 ;
        RECT 68.055 37.610 70.215 38.790 ;
        RECT 51.055 35.250 51.285 35.390 ;
        RECT 52.025 35.250 52.400 35.390 ;
        RECT 51.055 35.085 52.400 35.250 ;
        RECT 55.055 35.120 57.215 36.300 ;
        RECT 68.055 35.950 70.215 37.130 ;
        RECT 51.055 34.930 51.285 35.085 ;
        RECT 52.025 34.930 52.400 35.085 ;
        RECT 48.435 34.520 49.610 34.730 ;
        RECT 40.195 32.570 40.525 32.720 ;
        RECT 41.355 32.570 41.585 32.720 ;
        RECT 40.195 32.415 41.585 32.570 ;
        RECT 40.195 32.260 40.525 32.415 ;
        RECT 41.355 32.260 41.585 32.415 ;
        RECT 43.685 32.570 43.915 32.720 ;
        RECT 44.745 32.570 44.975 32.720 ;
        RECT 47.365 32.570 47.675 33.245 ;
        RECT 48.420 32.805 51.865 33.015 ;
        RECT 48.445 32.660 48.865 32.805 ;
        RECT 51.445 32.660 51.865 32.805 ;
        RECT 52.160 32.610 52.400 34.930 ;
        RECT 55.055 33.460 57.215 34.640 ;
        RECT 68.055 34.290 70.215 35.470 ;
        RECT 43.685 32.410 47.675 32.570 ;
        RECT 48.055 32.480 48.285 32.610 ;
        RECT 49.025 32.480 49.255 32.610 ;
        RECT 43.685 32.260 43.915 32.410 ;
        RECT 44.745 32.260 44.975 32.410 ;
        RECT 47.365 32.360 47.675 32.410 ;
        RECT 48.010 32.295 49.255 32.480 ;
        RECT 40.195 32.100 40.430 32.260 ;
        RECT 40.730 32.100 41.150 32.210 ;
        RECT 44.120 32.100 44.540 32.210 ;
        RECT 48.055 32.150 48.285 32.295 ;
        RECT 49.025 32.150 49.255 32.295 ;
        RECT 51.055 32.470 51.285 32.610 ;
        RECT 52.025 32.470 52.400 32.610 ;
        RECT 51.055 32.305 52.400 32.470 ;
        RECT 51.055 32.150 51.285 32.305 ;
        RECT 52.025 32.150 52.400 32.305 ;
        RECT 40.195 31.915 44.560 32.100 ;
        RECT 48.445 31.915 48.865 32.100 ;
        RECT 40.195 31.865 48.875 31.915 ;
        RECT 44.325 31.680 48.875 31.865 ;
        RECT 21.805 29.210 23.965 30.390 ;
        RECT 34.805 30.040 36.965 31.220 ;
        RECT 49.045 31.085 49.230 32.150 ;
        RECT 47.490 30.900 49.230 31.085 ;
        RECT 47.490 30.685 47.675 30.900 ;
        RECT 47.385 29.800 47.695 30.685 ;
        RECT 52.160 30.245 52.400 32.150 ;
        RECT 55.055 31.800 57.215 32.980 ;
        RECT 68.055 32.630 70.215 33.810 ;
        RECT 48.410 30.045 52.400 30.245 ;
        RECT 55.055 30.140 57.215 31.320 ;
        RECT 68.055 30.970 70.215 32.150 ;
        RECT 48.455 29.880 48.875 30.045 ;
        RECT 51.445 29.880 51.865 30.045 ;
        RECT 52.160 29.830 52.400 30.045 ;
        RECT 47.490 29.700 47.695 29.800 ;
        RECT 48.065 29.700 48.295 29.830 ;
        RECT 49.035 29.700 49.265 29.830 ;
        RECT 21.805 27.550 23.965 28.730 ;
        RECT 34.805 28.380 36.965 29.560 ;
        RECT 47.490 29.515 49.265 29.700 ;
        RECT 48.065 29.370 48.295 29.515 ;
        RECT 49.035 29.370 49.265 29.515 ;
        RECT 51.055 29.685 51.285 29.830 ;
        RECT 52.025 29.685 52.400 29.830 ;
        RECT 51.055 29.520 52.400 29.685 ;
        RECT 51.055 29.370 51.285 29.520 ;
        RECT 52.025 29.370 52.400 29.520 ;
        RECT 48.455 29.195 48.875 29.320 ;
        RECT 39.600 29.090 48.875 29.195 ;
        RECT 39.600 28.940 48.855 29.090 ;
        RECT 21.805 25.890 23.965 27.070 ;
        RECT 34.805 26.720 36.965 27.900 ;
        RECT 21.805 24.230 23.965 25.410 ;
        RECT 34.805 25.060 36.965 26.240 ;
        RECT 21.805 22.570 23.965 23.750 ;
        RECT 34.805 23.400 36.965 24.580 ;
        RECT 39.600 22.940 39.855 28.940 ;
        RECT 47.970 27.195 48.280 28.080 ;
        RECT 52.160 27.430 52.400 29.370 ;
        RECT 55.055 28.480 57.215 29.660 ;
        RECT 68.055 29.310 70.215 30.490 ;
        RECT 48.465 27.330 52.400 27.430 ;
        RECT 48.455 27.270 52.400 27.330 ;
        RECT 48.075 27.050 48.275 27.195 ;
        RECT 48.455 27.100 48.875 27.270 ;
        RECT 48.065 26.880 48.295 27.050 ;
        RECT 49.035 26.880 49.265 27.050 ;
        RECT 48.065 26.740 49.265 26.880 ;
        RECT 55.055 26.820 57.215 28.000 ;
        RECT 68.055 27.650 70.215 28.830 ;
        RECT 48.065 26.590 48.295 26.740 ;
        RECT 49.035 26.590 49.265 26.740 ;
        RECT 55.055 25.160 57.215 26.340 ;
        RECT 68.055 25.990 70.215 27.170 ;
        RECT 55.055 23.500 57.215 24.680 ;
        RECT 68.055 24.330 70.215 25.510 ;
        RECT 34.800 22.565 39.855 22.940 ;
        RECT 68.055 22.670 70.215 23.850 ;
      LAYER via ;
        RECT 44.495 77.965 44.755 78.225 ;
        RECT 44.495 77.645 44.755 77.905 ;
        RECT 44.000 74.605 44.260 74.865 ;
        RECT 43.955 71.720 44.215 71.980 ;
        RECT 43.955 71.400 44.215 71.660 ;
        RECT 46.390 67.025 46.650 67.285 ;
        RECT 45.290 66.325 45.550 66.585 ;
        RECT 47.040 66.335 47.300 66.595 ;
        RECT 46.380 64.685 46.640 64.945 ;
        RECT 48.160 64.685 48.420 64.945 ;
        RECT 44.000 63.965 44.260 64.225 ;
        RECT 45.290 63.975 45.550 64.235 ;
        RECT 47.050 62.685 47.310 62.945 ;
        RECT 48.200 62.685 48.460 62.945 ;
        RECT 42.930 60.815 43.190 61.075 ;
        RECT 42.930 60.495 43.190 60.755 ;
        RECT 42.930 60.175 43.190 60.435 ;
        RECT 48.030 60.355 48.290 60.615 ;
        RECT 48.030 60.035 48.290 60.295 ;
        RECT 48.030 59.715 48.290 59.975 ;
        RECT 46.270 54.520 46.530 54.780 ;
        RECT 46.590 54.520 46.850 54.780 ;
        RECT 45.320 50.135 45.580 50.395 ;
        RECT 45.320 49.815 45.580 50.075 ;
        RECT 45.320 49.495 45.580 49.755 ;
        RECT 45.320 46.070 45.580 46.330 ;
        RECT 45.320 45.750 45.580 46.010 ;
        RECT 45.320 45.430 45.580 45.690 ;
        RECT 45.320 43.050 45.580 43.310 ;
        RECT 45.320 42.730 45.580 42.990 ;
        RECT 45.320 42.410 45.580 42.670 ;
        RECT 45.320 39.890 45.580 40.150 ;
        RECT 45.320 39.570 45.580 39.830 ;
        RECT 45.320 39.250 45.580 39.510 ;
        RECT 45.320 36.735 45.580 36.995 ;
        RECT 45.320 36.415 45.580 36.675 ;
        RECT 45.320 36.095 45.580 36.355 ;
        RECT 46.290 35.025 46.550 35.285 ;
        RECT 46.610 35.025 46.870 35.285 ;
        RECT 47.390 32.830 47.650 33.090 ;
        RECT 47.390 32.510 47.650 32.770 ;
        RECT 47.410 30.270 47.670 30.530 ;
        RECT 47.410 29.950 47.670 30.210 ;
        RECT 47.995 27.665 48.255 27.925 ;
        RECT 47.995 27.345 48.255 27.605 ;
      LAYER met2 ;
        RECT 44.395 77.495 44.855 78.375 ;
        RECT 44.535 77.120 44.755 77.495 ;
        RECT 43.425 76.900 44.755 77.120 ;
        RECT 43.425 69.860 43.645 76.900 ;
        RECT 43.915 74.490 44.345 74.980 ;
        RECT 43.995 72.130 44.265 74.490 ;
        RECT 43.855 71.250 44.315 72.130 ;
        RECT 42.940 69.640 43.645 69.860 ;
        RECT 42.940 61.105 43.160 69.640 ;
        RECT 43.995 64.340 44.265 71.250 ;
        RECT 46.305 66.910 46.735 67.400 ;
        RECT 45.305 66.700 45.575 66.800 ;
        RECT 45.205 66.210 45.635 66.700 ;
        RECT 45.305 64.350 45.575 66.210 ;
        RECT 46.375 65.060 46.645 66.910 ;
        RECT 46.955 66.220 47.385 66.710 ;
        RECT 46.295 64.570 46.725 65.060 ;
        RECT 46.375 64.500 46.645 64.570 ;
        RECT 43.915 63.850 44.345 64.340 ;
        RECT 45.205 63.860 45.635 64.350 ;
        RECT 47.025 63.060 47.305 66.220 ;
        RECT 48.075 64.570 48.505 65.060 ;
        RECT 48.185 63.060 48.455 64.570 ;
        RECT 46.965 62.570 47.395 63.060 ;
        RECT 48.115 62.570 48.545 63.060 ;
        RECT 48.175 61.315 48.480 62.570 ;
        RECT 42.815 60.150 43.305 61.105 ;
        RECT 47.385 61.010 48.480 61.315 ;
        RECT 46.095 54.510 47.020 54.795 ;
        RECT 44.795 53.925 45.970 54.415 ;
        RECT 45.170 50.470 45.720 53.925 ;
        RECT 45.170 50.410 45.725 50.470 ;
        RECT 45.175 49.420 45.725 50.410 ;
        RECT 44.795 48.595 45.970 49.085 ;
        RECT 45.175 46.405 45.720 48.595 ;
        RECT 45.175 45.355 45.725 46.405 ;
        RECT 44.795 43.265 45.970 43.755 ;
        RECT 45.175 42.335 45.725 43.265 ;
        RECT 45.175 39.255 45.725 40.225 ;
        RECT 45.170 39.175 45.725 39.255 ;
        RECT 45.170 38.425 45.720 39.175 ;
        RECT 44.795 37.935 45.970 38.425 ;
        RECT 45.175 36.020 45.725 37.070 ;
        RECT 45.190 33.095 45.715 36.020 ;
        RECT 46.500 35.300 46.705 54.510 ;
        RECT 46.115 35.015 47.040 35.300 ;
        RECT 47.385 33.195 47.690 61.010 ;
        RECT 47.950 59.700 48.370 60.635 ;
        RECT 47.950 59.650 48.280 59.700 ;
        RECT 44.795 32.605 45.970 33.095 ;
        RECT 47.315 32.410 47.725 33.195 ;
        RECT 47.385 30.635 47.690 32.410 ;
        RECT 47.335 29.850 47.745 30.635 ;
        RECT 47.385 29.660 47.690 29.850 ;
        RECT 48.055 28.030 48.280 59.650 ;
        RECT 47.920 27.245 48.330 28.030 ;
      LAYER via2 ;
        RECT 45.045 54.030 45.325 54.310 ;
        RECT 45.445 54.030 45.725 54.310 ;
        RECT 45.045 48.700 45.325 48.980 ;
        RECT 45.445 48.700 45.725 48.980 ;
        RECT 45.045 43.370 45.325 43.650 ;
        RECT 45.445 43.370 45.725 43.650 ;
        RECT 45.045 38.040 45.325 38.320 ;
        RECT 45.445 38.040 45.725 38.320 ;
        RECT 45.045 32.710 45.325 32.990 ;
        RECT 45.445 32.710 45.725 32.990 ;
      LAYER met3 ;
        RECT 44.820 53.875 45.945 54.465 ;
        RECT 44.820 48.545 45.945 49.135 ;
        RECT 44.820 43.215 45.945 43.805 ;
        RECT 44.820 37.885 45.945 38.475 ;
        RECT 44.820 32.555 45.945 33.145 ;
      LAYER via3 ;
        RECT 45.025 54.010 45.345 54.330 ;
        RECT 45.425 54.010 45.745 54.330 ;
        RECT 45.025 48.680 45.345 49.000 ;
        RECT 45.425 48.680 45.745 49.000 ;
        RECT 45.025 43.350 45.345 43.670 ;
        RECT 45.425 43.350 45.745 43.670 ;
        RECT 45.025 38.020 45.345 38.340 ;
        RECT 45.425 38.020 45.745 38.340 ;
        RECT 45.025 32.690 45.345 33.010 ;
        RECT 45.425 32.690 45.745 33.010 ;
      LAYER met4 ;
        RECT 44.815 54.415 45.955 54.470 ;
        RECT 47.145 54.415 52.755 55.485 ;
        RECT 44.815 53.925 52.755 54.415 ;
        RECT 44.815 53.870 45.955 53.925 ;
        RECT 47.145 52.875 52.755 53.925 ;
        RECT 44.815 49.085 45.955 49.140 ;
        RECT 47.145 49.085 52.755 50.155 ;
        RECT 44.815 48.595 52.755 49.085 ;
        RECT 44.815 48.540 45.955 48.595 ;
        RECT 47.145 47.545 52.755 48.595 ;
        RECT 44.815 43.755 45.955 43.810 ;
        RECT 47.145 43.755 52.755 44.825 ;
        RECT 44.815 43.265 52.755 43.755 ;
        RECT 44.815 43.210 45.955 43.265 ;
        RECT 47.145 42.215 52.755 43.265 ;
        RECT 44.815 38.425 45.955 38.480 ;
        RECT 47.150 38.425 52.760 39.495 ;
        RECT 44.815 37.935 52.760 38.425 ;
        RECT 44.815 37.880 45.955 37.935 ;
        RECT 47.150 36.885 52.760 37.935 ;
        RECT 44.815 33.095 45.955 33.150 ;
        RECT 47.150 33.095 52.760 34.165 ;
        RECT 44.815 32.605 52.760 33.095 ;
        RECT 44.815 32.550 45.955 32.605 ;
        RECT 47.150 31.555 52.760 32.605 ;
  END
END sky130_ef_ip__rc_osc_500k_DI
END LIBRARY


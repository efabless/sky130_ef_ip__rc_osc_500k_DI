magic
tech sky130A
magscale 1 2
timestamp 1528473026
<< checkpaint >>
rect -1140 -1260 12104 30103
<< via1 >>
rect 3735 18647 3787 18699
rect 3799 18647 3851 18699
rect 3863 18647 3915 18699
rect 3927 18647 3979 18699
rect 4103 18647 4155 18699
rect 4167 18647 4219 18699
rect 4231 18647 4283 18699
rect 4409 18646 4461 18698
rect 6469 18647 6521 18699
rect 6533 18647 6585 18699
rect 6597 18647 6649 18699
rect 6661 18647 6713 18699
rect 6837 18647 6889 18699
rect 6901 18647 6953 18699
rect 6965 18647 7017 18699
rect 7143 18646 7195 18698
rect 3735 18557 3787 18609
rect 3799 18557 3851 18609
rect 3863 18557 3915 18609
rect 3927 18557 3979 18609
rect 4103 18557 4155 18609
rect 4167 18557 4219 18609
rect 4231 18557 4283 18609
rect 4409 18556 4461 18608
rect 6469 18557 6521 18609
rect 6533 18557 6585 18609
rect 6597 18557 6649 18609
rect 6661 18557 6713 18609
rect 6837 18557 6889 18609
rect 6901 18557 6953 18609
rect 6965 18557 7017 18609
rect 7143 18556 7195 18608
<< metal2 >>
rect 5289 27537 5401 28843
rect 5933 27643 6045 28843
rect 5147 27509 5401 27537
rect 3723 18699 4480 18706
rect 3723 18647 3735 18699
rect 3787 18697 3799 18699
rect 3851 18697 3863 18699
rect 3915 18697 3927 18699
rect 3979 18697 4103 18699
rect 4155 18697 4167 18699
rect 4219 18697 4231 18699
rect 4283 18698 4480 18699
rect 4283 18697 4409 18698
rect 3794 18647 3799 18697
rect 4034 18647 4103 18697
rect 4160 18647 4167 18697
rect 3723 18641 3738 18647
rect 3794 18641 3818 18647
rect 3874 18641 3898 18647
rect 3954 18641 3978 18647
rect 4034 18641 4104 18647
rect 4160 18641 4184 18647
rect 4240 18641 4264 18647
rect 4320 18641 4344 18697
rect 4400 18646 4409 18697
rect 4461 18646 4480 18698
rect 4400 18641 4480 18646
rect 3723 18609 4480 18641
rect 3723 18557 3735 18609
rect 3787 18578 3799 18609
rect 3851 18578 3863 18609
rect 3915 18578 3927 18609
rect 3979 18578 4103 18609
rect 4155 18578 4167 18609
rect 4219 18578 4231 18609
rect 4283 18608 4480 18609
rect 4283 18578 4409 18608
rect 3794 18557 3799 18578
rect 4034 18557 4103 18578
rect 4160 18557 4167 18578
rect 3723 18522 3738 18557
rect 3794 18522 3818 18557
rect 3874 18522 3898 18557
rect 3954 18522 3978 18557
rect 4034 18522 4104 18557
rect 4160 18522 4184 18557
rect 4240 18522 4264 18557
rect 4320 18522 4344 18578
rect 4400 18556 4409 18578
rect 4461 18556 4480 18608
rect 5147 18580 5175 27509
rect 5289 27403 5401 27509
rect 5924 27403 6045 27643
rect 5924 27401 5952 27403
rect 5883 27373 5952 27401
rect 5883 18580 5911 27373
rect 6453 18699 7210 18706
rect 6453 18697 6469 18699
rect 6521 18697 6533 18699
rect 6585 18697 6597 18699
rect 6649 18697 6661 18699
rect 6713 18697 6837 18699
rect 6889 18697 6901 18699
rect 6953 18697 6965 18699
rect 7017 18698 7210 18699
rect 7017 18697 7143 18698
rect 6453 18641 6468 18697
rect 6524 18647 6533 18697
rect 6524 18641 6548 18647
rect 6604 18641 6628 18647
rect 6684 18641 6708 18647
rect 6764 18641 6834 18697
rect 6890 18647 6901 18697
rect 6890 18641 6914 18647
rect 6970 18641 6994 18647
rect 7050 18641 7074 18697
rect 7130 18646 7143 18697
rect 7195 18646 7210 18698
rect 7130 18641 7210 18646
rect 6453 18609 7210 18641
rect 4400 18522 4480 18556
rect 3723 18506 4480 18522
rect 6453 18578 6469 18609
rect 6521 18578 6533 18609
rect 6585 18578 6597 18609
rect 6649 18578 6661 18609
rect 6713 18578 6837 18609
rect 6889 18578 6901 18609
rect 6953 18578 6965 18609
rect 7017 18608 7210 18609
rect 7017 18578 7143 18608
rect 6453 18522 6468 18578
rect 6524 18557 6533 18578
rect 6524 18522 6548 18557
rect 6604 18522 6628 18557
rect 6684 18522 6708 18557
rect 6764 18522 6834 18578
rect 6890 18557 6901 18578
rect 6890 18522 6914 18557
rect 6970 18522 6994 18557
rect 7050 18522 7074 18578
rect 7130 18556 7143 18578
rect 7195 18556 7210 18608
rect 7130 18522 7210 18556
rect 6453 18506 7210 18522
<< via2 >>
rect 3738 18647 3787 18697
rect 3787 18647 3794 18697
rect 3818 18647 3851 18697
rect 3851 18647 3863 18697
rect 3863 18647 3874 18697
rect 3898 18647 3915 18697
rect 3915 18647 3927 18697
rect 3927 18647 3954 18697
rect 3978 18647 3979 18697
rect 3979 18647 4034 18697
rect 4104 18647 4155 18697
rect 4155 18647 4160 18697
rect 4184 18647 4219 18697
rect 4219 18647 4231 18697
rect 4231 18647 4240 18697
rect 4264 18647 4283 18697
rect 4283 18647 4320 18697
rect 3738 18641 3794 18647
rect 3818 18641 3874 18647
rect 3898 18641 3954 18647
rect 3978 18641 4034 18647
rect 4104 18641 4160 18647
rect 4184 18641 4240 18647
rect 4264 18641 4320 18647
rect 4344 18641 4400 18697
rect 3738 18557 3787 18578
rect 3787 18557 3794 18578
rect 3818 18557 3851 18578
rect 3851 18557 3863 18578
rect 3863 18557 3874 18578
rect 3898 18557 3915 18578
rect 3915 18557 3927 18578
rect 3927 18557 3954 18578
rect 3978 18557 3979 18578
rect 3979 18557 4034 18578
rect 4104 18557 4155 18578
rect 4155 18557 4160 18578
rect 4184 18557 4219 18578
rect 4219 18557 4231 18578
rect 4231 18557 4240 18578
rect 4264 18557 4283 18578
rect 4283 18557 4320 18578
rect 3738 18522 3794 18557
rect 3818 18522 3874 18557
rect 3898 18522 3954 18557
rect 3978 18522 4034 18557
rect 4104 18522 4160 18557
rect 4184 18522 4240 18557
rect 4264 18522 4320 18557
rect 4344 18522 4400 18578
rect 6468 18647 6469 18697
rect 6469 18647 6521 18697
rect 6521 18647 6524 18697
rect 6548 18647 6585 18697
rect 6585 18647 6597 18697
rect 6597 18647 6604 18697
rect 6628 18647 6649 18697
rect 6649 18647 6661 18697
rect 6661 18647 6684 18697
rect 6708 18647 6713 18697
rect 6713 18647 6764 18697
rect 6468 18641 6524 18647
rect 6548 18641 6604 18647
rect 6628 18641 6684 18647
rect 6708 18641 6764 18647
rect 6834 18647 6837 18697
rect 6837 18647 6889 18697
rect 6889 18647 6890 18697
rect 6914 18647 6953 18697
rect 6953 18647 6965 18697
rect 6965 18647 6970 18697
rect 6994 18647 7017 18697
rect 7017 18647 7050 18697
rect 6834 18641 6890 18647
rect 6914 18641 6970 18647
rect 6994 18641 7050 18647
rect 7074 18641 7130 18697
rect 6468 18557 6469 18578
rect 6469 18557 6521 18578
rect 6521 18557 6524 18578
rect 6548 18557 6585 18578
rect 6585 18557 6597 18578
rect 6597 18557 6604 18578
rect 6628 18557 6649 18578
rect 6649 18557 6661 18578
rect 6661 18557 6684 18578
rect 6708 18557 6713 18578
rect 6713 18557 6764 18578
rect 6468 18522 6524 18557
rect 6548 18522 6604 18557
rect 6628 18522 6684 18557
rect 6708 18522 6764 18557
rect 6834 18557 6837 18578
rect 6837 18557 6889 18578
rect 6889 18557 6890 18578
rect 6914 18557 6953 18578
rect 6953 18557 6965 18578
rect 6965 18557 6970 18578
rect 6994 18557 7017 18578
rect 7017 18557 7050 18578
rect 6834 18522 6890 18557
rect 6914 18522 6970 18557
rect 6994 18522 7050 18557
rect 7074 18522 7130 18578
rect 1714 18411 1770 18467
rect 1794 18411 1850 18467
rect 1874 18411 1930 18467
rect 1954 18411 2010 18467
rect 2380 18411 2436 18467
rect 2460 18411 2516 18467
rect 2540 18411 2596 18467
rect 2620 18411 2676 18467
rect 8428 18438 8484 18494
rect 8508 18438 8564 18494
rect 8588 18438 8644 18494
rect 8668 18438 8724 18494
rect 9094 18438 9150 18494
rect 9174 18438 9230 18494
rect 9254 18438 9310 18494
rect 9334 18438 9390 18494
rect 1714 18292 1770 18348
rect 1794 18292 1850 18348
rect 1874 18292 1930 18348
rect 1954 18292 2010 18348
rect 2380 18292 2436 18348
rect 2460 18292 2516 18348
rect 2540 18292 2596 18348
rect 2620 18292 2676 18348
rect 8428 18319 8484 18375
rect 8508 18319 8564 18375
rect 8588 18319 8644 18375
rect 8668 18319 8724 18375
rect 9094 18319 9150 18375
rect 9174 18319 9230 18375
rect 9254 18319 9310 18375
rect 9334 18319 9390 18375
rect 1714 6591 1770 6647
rect 1794 6591 1850 6647
rect 1874 6591 1930 6647
rect 1954 6591 2010 6647
rect 2380 6591 2436 6647
rect 2460 6591 2516 6647
rect 2540 6591 2596 6647
rect 2620 6591 2676 6647
rect 8428 6598 8484 6654
rect 8508 6598 8564 6654
rect 8588 6598 8644 6654
rect 8668 6598 8724 6654
rect 9094 6598 9150 6654
rect 9174 6598 9230 6654
rect 9254 6598 9310 6654
rect 9334 6598 9390 6654
rect 1714 6472 1770 6528
rect 1794 6472 1850 6528
rect 1874 6472 1930 6528
rect 1954 6472 2010 6528
rect 2380 6472 2436 6528
rect 2460 6472 2516 6528
rect 2540 6472 2596 6528
rect 2620 6472 2676 6528
rect 8428 6479 8484 6535
rect 8508 6479 8564 6535
rect 8588 6479 8644 6535
rect 8668 6479 8724 6535
rect 9094 6479 9150 6535
rect 9174 6479 9230 6535
rect 9254 6479 9310 6535
rect 9334 6479 9390 6535
<< metal3 >>
rect 3723 18701 4480 18706
rect 3723 18637 3734 18701
rect 3798 18637 3814 18701
rect 3878 18637 3894 18701
rect 3958 18637 3974 18701
rect 4038 18637 4100 18701
rect 4164 18637 4180 18701
rect 4244 18637 4260 18701
rect 4324 18697 4480 18701
rect 4324 18641 4344 18697
rect 4400 18641 4480 18697
rect 4324 18637 4480 18641
rect 1699 18471 2699 18625
rect 3723 18582 4480 18637
rect 3723 18518 3734 18582
rect 3798 18518 3814 18582
rect 3878 18518 3894 18582
rect 3958 18518 3974 18582
rect 4038 18518 4100 18582
rect 4164 18518 4180 18582
rect 4244 18518 4260 18582
rect 4324 18578 4480 18582
rect 4324 18522 4344 18578
rect 4400 18522 4480 18578
rect 4324 18518 4480 18522
rect 3723 18506 4480 18518
rect 6453 18701 7210 18706
rect 6453 18637 6464 18701
rect 6528 18637 6544 18701
rect 6608 18637 6624 18701
rect 6688 18637 6704 18701
rect 6768 18637 6830 18701
rect 6894 18637 6910 18701
rect 6974 18637 6990 18701
rect 7054 18697 7210 18701
rect 7054 18641 7074 18697
rect 7130 18641 7210 18697
rect 7054 18637 7210 18641
rect 6453 18582 7210 18637
rect 6453 18518 6464 18582
rect 6528 18518 6544 18582
rect 6608 18518 6624 18582
rect 6688 18518 6704 18582
rect 6768 18518 6830 18582
rect 6894 18518 6910 18582
rect 6974 18518 6990 18582
rect 7054 18578 7210 18582
rect 7054 18522 7074 18578
rect 7130 18522 7210 18578
rect 7054 18518 7210 18522
rect 6453 18506 7210 18518
rect 1699 18407 1710 18471
rect 1774 18407 1790 18471
rect 1854 18407 1870 18471
rect 1934 18407 1950 18471
rect 2014 18407 2376 18471
rect 2440 18407 2456 18471
rect 2520 18407 2536 18471
rect 2600 18407 2616 18471
rect 2680 18407 2699 18471
rect 1699 18352 2699 18407
rect 1699 18288 1710 18352
rect 1774 18288 1790 18352
rect 1854 18288 1870 18352
rect 1934 18288 1950 18352
rect 2014 18288 2376 18352
rect 2440 18288 2456 18352
rect 2520 18288 2536 18352
rect 2600 18288 2616 18352
rect 2680 18288 2699 18352
rect 8413 18498 9413 18645
rect 8413 18434 8424 18498
rect 8488 18434 8504 18498
rect 8568 18434 8584 18498
rect 8648 18434 8664 18498
rect 8728 18434 9090 18498
rect 9154 18434 9170 18498
rect 9234 18434 9250 18498
rect 9314 18434 9330 18498
rect 9394 18434 9413 18498
rect 8413 18379 9413 18434
rect 8413 18315 8424 18379
rect 8488 18315 8504 18379
rect 8568 18315 8584 18379
rect 8648 18315 8664 18379
rect 8728 18315 9090 18379
rect 9154 18315 9170 18379
rect 9234 18315 9250 18379
rect 9314 18315 9330 18379
rect 9394 18315 9413 18379
rect 8413 18303 9413 18315
rect 1699 18283 2699 18288
rect 1699 6651 2699 6805
rect 1699 6587 1710 6651
rect 1774 6587 1790 6651
rect 1854 6587 1870 6651
rect 1934 6587 1950 6651
rect 2014 6587 2376 6651
rect 2440 6587 2456 6651
rect 2520 6587 2536 6651
rect 2600 6587 2616 6651
rect 2680 6587 2699 6651
rect 1699 6532 2699 6587
rect 1699 6468 1710 6532
rect 1774 6468 1790 6532
rect 1854 6468 1870 6532
rect 1934 6468 1950 6532
rect 2014 6468 2376 6532
rect 2440 6468 2456 6532
rect 2520 6468 2536 6532
rect 2600 6468 2616 6532
rect 2680 6468 2699 6532
rect 1699 6463 2699 6468
rect 8413 6658 9413 6805
rect 8413 6594 8424 6658
rect 8488 6594 8504 6658
rect 8568 6594 8584 6658
rect 8648 6594 8664 6658
rect 8728 6594 9090 6658
rect 9154 6594 9170 6658
rect 9234 6594 9250 6658
rect 9314 6594 9330 6658
rect 9394 6594 9413 6658
rect 8413 6539 9413 6594
rect 8413 6475 8424 6539
rect 8488 6475 8504 6539
rect 8568 6475 8584 6539
rect 8648 6475 8664 6539
rect 8728 6475 9090 6539
rect 9154 6475 9170 6539
rect 9234 6475 9250 6539
rect 9314 6475 9330 6539
rect 9394 6475 9413 6539
rect 8413 6463 9413 6475
<< via3 >>
rect 3734 18697 3798 18701
rect 3734 18641 3738 18697
rect 3738 18641 3794 18697
rect 3794 18641 3798 18697
rect 3734 18637 3798 18641
rect 3814 18697 3878 18701
rect 3814 18641 3818 18697
rect 3818 18641 3874 18697
rect 3874 18641 3878 18697
rect 3814 18637 3878 18641
rect 3894 18697 3958 18701
rect 3894 18641 3898 18697
rect 3898 18641 3954 18697
rect 3954 18641 3958 18697
rect 3894 18637 3958 18641
rect 3974 18697 4038 18701
rect 3974 18641 3978 18697
rect 3978 18641 4034 18697
rect 4034 18641 4038 18697
rect 3974 18637 4038 18641
rect 4100 18697 4164 18701
rect 4100 18641 4104 18697
rect 4104 18641 4160 18697
rect 4160 18641 4164 18697
rect 4100 18637 4164 18641
rect 4180 18697 4244 18701
rect 4180 18641 4184 18697
rect 4184 18641 4240 18697
rect 4240 18641 4244 18697
rect 4180 18637 4244 18641
rect 4260 18697 4324 18701
rect 4260 18641 4264 18697
rect 4264 18641 4320 18697
rect 4320 18641 4324 18697
rect 4260 18637 4324 18641
rect 3734 18578 3798 18582
rect 3734 18522 3738 18578
rect 3738 18522 3794 18578
rect 3794 18522 3798 18578
rect 3734 18518 3798 18522
rect 3814 18578 3878 18582
rect 3814 18522 3818 18578
rect 3818 18522 3874 18578
rect 3874 18522 3878 18578
rect 3814 18518 3878 18522
rect 3894 18578 3958 18582
rect 3894 18522 3898 18578
rect 3898 18522 3954 18578
rect 3954 18522 3958 18578
rect 3894 18518 3958 18522
rect 3974 18578 4038 18582
rect 3974 18522 3978 18578
rect 3978 18522 4034 18578
rect 4034 18522 4038 18578
rect 3974 18518 4038 18522
rect 4100 18578 4164 18582
rect 4100 18522 4104 18578
rect 4104 18522 4160 18578
rect 4160 18522 4164 18578
rect 4100 18518 4164 18522
rect 4180 18578 4244 18582
rect 4180 18522 4184 18578
rect 4184 18522 4240 18578
rect 4240 18522 4244 18578
rect 4180 18518 4244 18522
rect 4260 18578 4324 18582
rect 4260 18522 4264 18578
rect 4264 18522 4320 18578
rect 4320 18522 4324 18578
rect 4260 18518 4324 18522
rect 6464 18697 6528 18701
rect 6464 18641 6468 18697
rect 6468 18641 6524 18697
rect 6524 18641 6528 18697
rect 6464 18637 6528 18641
rect 6544 18697 6608 18701
rect 6544 18641 6548 18697
rect 6548 18641 6604 18697
rect 6604 18641 6608 18697
rect 6544 18637 6608 18641
rect 6624 18697 6688 18701
rect 6624 18641 6628 18697
rect 6628 18641 6684 18697
rect 6684 18641 6688 18697
rect 6624 18637 6688 18641
rect 6704 18697 6768 18701
rect 6704 18641 6708 18697
rect 6708 18641 6764 18697
rect 6764 18641 6768 18697
rect 6704 18637 6768 18641
rect 6830 18697 6894 18701
rect 6830 18641 6834 18697
rect 6834 18641 6890 18697
rect 6890 18641 6894 18697
rect 6830 18637 6894 18641
rect 6910 18697 6974 18701
rect 6910 18641 6914 18697
rect 6914 18641 6970 18697
rect 6970 18641 6974 18697
rect 6910 18637 6974 18641
rect 6990 18697 7054 18701
rect 6990 18641 6994 18697
rect 6994 18641 7050 18697
rect 7050 18641 7054 18697
rect 6990 18637 7054 18641
rect 6464 18578 6528 18582
rect 6464 18522 6468 18578
rect 6468 18522 6524 18578
rect 6524 18522 6528 18578
rect 6464 18518 6528 18522
rect 6544 18578 6608 18582
rect 6544 18522 6548 18578
rect 6548 18522 6604 18578
rect 6604 18522 6608 18578
rect 6544 18518 6608 18522
rect 6624 18578 6688 18582
rect 6624 18522 6628 18578
rect 6628 18522 6684 18578
rect 6684 18522 6688 18578
rect 6624 18518 6688 18522
rect 6704 18578 6768 18582
rect 6704 18522 6708 18578
rect 6708 18522 6764 18578
rect 6764 18522 6768 18578
rect 6704 18518 6768 18522
rect 6830 18578 6894 18582
rect 6830 18522 6834 18578
rect 6834 18522 6890 18578
rect 6890 18522 6894 18578
rect 6830 18518 6894 18522
rect 6910 18578 6974 18582
rect 6910 18522 6914 18578
rect 6914 18522 6970 18578
rect 6970 18522 6974 18578
rect 6910 18518 6974 18522
rect 6990 18578 7054 18582
rect 6990 18522 6994 18578
rect 6994 18522 7050 18578
rect 7050 18522 7054 18578
rect 6990 18518 7054 18522
rect 1710 18467 1774 18471
rect 1710 18411 1714 18467
rect 1714 18411 1770 18467
rect 1770 18411 1774 18467
rect 1710 18407 1774 18411
rect 1790 18467 1854 18471
rect 1790 18411 1794 18467
rect 1794 18411 1850 18467
rect 1850 18411 1854 18467
rect 1790 18407 1854 18411
rect 1870 18467 1934 18471
rect 1870 18411 1874 18467
rect 1874 18411 1930 18467
rect 1930 18411 1934 18467
rect 1870 18407 1934 18411
rect 1950 18467 2014 18471
rect 1950 18411 1954 18467
rect 1954 18411 2010 18467
rect 2010 18411 2014 18467
rect 1950 18407 2014 18411
rect 2376 18467 2440 18471
rect 2376 18411 2380 18467
rect 2380 18411 2436 18467
rect 2436 18411 2440 18467
rect 2376 18407 2440 18411
rect 2456 18467 2520 18471
rect 2456 18411 2460 18467
rect 2460 18411 2516 18467
rect 2516 18411 2520 18467
rect 2456 18407 2520 18411
rect 2536 18467 2600 18471
rect 2536 18411 2540 18467
rect 2540 18411 2596 18467
rect 2596 18411 2600 18467
rect 2536 18407 2600 18411
rect 2616 18467 2680 18471
rect 2616 18411 2620 18467
rect 2620 18411 2676 18467
rect 2676 18411 2680 18467
rect 2616 18407 2680 18411
rect 1710 18348 1774 18352
rect 1710 18292 1714 18348
rect 1714 18292 1770 18348
rect 1770 18292 1774 18348
rect 1710 18288 1774 18292
rect 1790 18348 1854 18352
rect 1790 18292 1794 18348
rect 1794 18292 1850 18348
rect 1850 18292 1854 18348
rect 1790 18288 1854 18292
rect 1870 18348 1934 18352
rect 1870 18292 1874 18348
rect 1874 18292 1930 18348
rect 1930 18292 1934 18348
rect 1870 18288 1934 18292
rect 1950 18348 2014 18352
rect 1950 18292 1954 18348
rect 1954 18292 2010 18348
rect 2010 18292 2014 18348
rect 1950 18288 2014 18292
rect 2376 18348 2440 18352
rect 2376 18292 2380 18348
rect 2380 18292 2436 18348
rect 2436 18292 2440 18348
rect 2376 18288 2440 18292
rect 2456 18348 2520 18352
rect 2456 18292 2460 18348
rect 2460 18292 2516 18348
rect 2516 18292 2520 18348
rect 2456 18288 2520 18292
rect 2536 18348 2600 18352
rect 2536 18292 2540 18348
rect 2540 18292 2596 18348
rect 2596 18292 2600 18348
rect 2536 18288 2600 18292
rect 2616 18348 2680 18352
rect 2616 18292 2620 18348
rect 2620 18292 2676 18348
rect 2676 18292 2680 18348
rect 2616 18288 2680 18292
rect 8424 18494 8488 18498
rect 8424 18438 8428 18494
rect 8428 18438 8484 18494
rect 8484 18438 8488 18494
rect 8424 18434 8488 18438
rect 8504 18494 8568 18498
rect 8504 18438 8508 18494
rect 8508 18438 8564 18494
rect 8564 18438 8568 18494
rect 8504 18434 8568 18438
rect 8584 18494 8648 18498
rect 8584 18438 8588 18494
rect 8588 18438 8644 18494
rect 8644 18438 8648 18494
rect 8584 18434 8648 18438
rect 8664 18494 8728 18498
rect 8664 18438 8668 18494
rect 8668 18438 8724 18494
rect 8724 18438 8728 18494
rect 8664 18434 8728 18438
rect 9090 18494 9154 18498
rect 9090 18438 9094 18494
rect 9094 18438 9150 18494
rect 9150 18438 9154 18494
rect 9090 18434 9154 18438
rect 9170 18494 9234 18498
rect 9170 18438 9174 18494
rect 9174 18438 9230 18494
rect 9230 18438 9234 18494
rect 9170 18434 9234 18438
rect 9250 18494 9314 18498
rect 9250 18438 9254 18494
rect 9254 18438 9310 18494
rect 9310 18438 9314 18494
rect 9250 18434 9314 18438
rect 9330 18494 9394 18498
rect 9330 18438 9334 18494
rect 9334 18438 9390 18494
rect 9390 18438 9394 18494
rect 9330 18434 9394 18438
rect 8424 18375 8488 18379
rect 8424 18319 8428 18375
rect 8428 18319 8484 18375
rect 8484 18319 8488 18375
rect 8424 18315 8488 18319
rect 8504 18375 8568 18379
rect 8504 18319 8508 18375
rect 8508 18319 8564 18375
rect 8564 18319 8568 18375
rect 8504 18315 8568 18319
rect 8584 18375 8648 18379
rect 8584 18319 8588 18375
rect 8588 18319 8644 18375
rect 8644 18319 8648 18375
rect 8584 18315 8648 18319
rect 8664 18375 8728 18379
rect 8664 18319 8668 18375
rect 8668 18319 8724 18375
rect 8724 18319 8728 18375
rect 8664 18315 8728 18319
rect 9090 18375 9154 18379
rect 9090 18319 9094 18375
rect 9094 18319 9150 18375
rect 9150 18319 9154 18375
rect 9090 18315 9154 18319
rect 9170 18375 9234 18379
rect 9170 18319 9174 18375
rect 9174 18319 9230 18375
rect 9230 18319 9234 18375
rect 9170 18315 9234 18319
rect 9250 18375 9314 18379
rect 9250 18319 9254 18375
rect 9254 18319 9310 18375
rect 9310 18319 9314 18375
rect 9250 18315 9314 18319
rect 9330 18375 9394 18379
rect 9330 18319 9334 18375
rect 9334 18319 9390 18375
rect 9390 18319 9394 18375
rect 9330 18315 9394 18319
rect 1710 6647 1774 6651
rect 1710 6591 1714 6647
rect 1714 6591 1770 6647
rect 1770 6591 1774 6647
rect 1710 6587 1774 6591
rect 1790 6647 1854 6651
rect 1790 6591 1794 6647
rect 1794 6591 1850 6647
rect 1850 6591 1854 6647
rect 1790 6587 1854 6591
rect 1870 6647 1934 6651
rect 1870 6591 1874 6647
rect 1874 6591 1930 6647
rect 1930 6591 1934 6647
rect 1870 6587 1934 6591
rect 1950 6647 2014 6651
rect 1950 6591 1954 6647
rect 1954 6591 2010 6647
rect 2010 6591 2014 6647
rect 1950 6587 2014 6591
rect 2376 6647 2440 6651
rect 2376 6591 2380 6647
rect 2380 6591 2436 6647
rect 2436 6591 2440 6647
rect 2376 6587 2440 6591
rect 2456 6647 2520 6651
rect 2456 6591 2460 6647
rect 2460 6591 2516 6647
rect 2516 6591 2520 6647
rect 2456 6587 2520 6591
rect 2536 6647 2600 6651
rect 2536 6591 2540 6647
rect 2540 6591 2596 6647
rect 2596 6591 2600 6647
rect 2536 6587 2600 6591
rect 2616 6647 2680 6651
rect 2616 6591 2620 6647
rect 2620 6591 2676 6647
rect 2676 6591 2680 6647
rect 2616 6587 2680 6591
rect 1710 6528 1774 6532
rect 1710 6472 1714 6528
rect 1714 6472 1770 6528
rect 1770 6472 1774 6528
rect 1710 6468 1774 6472
rect 1790 6528 1854 6532
rect 1790 6472 1794 6528
rect 1794 6472 1850 6528
rect 1850 6472 1854 6528
rect 1790 6468 1854 6472
rect 1870 6528 1934 6532
rect 1870 6472 1874 6528
rect 1874 6472 1930 6528
rect 1930 6472 1934 6528
rect 1870 6468 1934 6472
rect 1950 6528 2014 6532
rect 1950 6472 1954 6528
rect 1954 6472 2010 6528
rect 2010 6472 2014 6528
rect 1950 6468 2014 6472
rect 2376 6528 2440 6532
rect 2376 6472 2380 6528
rect 2380 6472 2436 6528
rect 2436 6472 2440 6528
rect 2376 6468 2440 6472
rect 2456 6528 2520 6532
rect 2456 6472 2460 6528
rect 2460 6472 2516 6528
rect 2516 6472 2520 6528
rect 2456 6468 2520 6472
rect 2536 6528 2600 6532
rect 2536 6472 2540 6528
rect 2540 6472 2596 6528
rect 2596 6472 2600 6528
rect 2536 6468 2600 6472
rect 2616 6528 2680 6532
rect 2616 6472 2620 6528
rect 2620 6472 2676 6528
rect 2676 6472 2680 6528
rect 2616 6468 2680 6472
rect 8424 6654 8488 6658
rect 8424 6598 8428 6654
rect 8428 6598 8484 6654
rect 8484 6598 8488 6654
rect 8424 6594 8488 6598
rect 8504 6654 8568 6658
rect 8504 6598 8508 6654
rect 8508 6598 8564 6654
rect 8564 6598 8568 6654
rect 8504 6594 8568 6598
rect 8584 6654 8648 6658
rect 8584 6598 8588 6654
rect 8588 6598 8644 6654
rect 8644 6598 8648 6654
rect 8584 6594 8648 6598
rect 8664 6654 8728 6658
rect 8664 6598 8668 6654
rect 8668 6598 8724 6654
rect 8724 6598 8728 6654
rect 8664 6594 8728 6598
rect 9090 6654 9154 6658
rect 9090 6598 9094 6654
rect 9094 6598 9150 6654
rect 9150 6598 9154 6654
rect 9090 6594 9154 6598
rect 9170 6654 9234 6658
rect 9170 6598 9174 6654
rect 9174 6598 9230 6654
rect 9230 6598 9234 6654
rect 9170 6594 9234 6598
rect 9250 6654 9314 6658
rect 9250 6598 9254 6654
rect 9254 6598 9310 6654
rect 9310 6598 9314 6654
rect 9250 6594 9314 6598
rect 9330 6654 9394 6658
rect 9330 6598 9334 6654
rect 9334 6598 9390 6654
rect 9390 6598 9394 6654
rect 9330 6594 9394 6598
rect 8424 6535 8488 6539
rect 8424 6479 8428 6535
rect 8428 6479 8484 6535
rect 8484 6479 8488 6535
rect 8424 6475 8488 6479
rect 8504 6535 8568 6539
rect 8504 6479 8508 6535
rect 8508 6479 8564 6535
rect 8564 6479 8568 6535
rect 8504 6475 8568 6479
rect 8584 6535 8648 6539
rect 8584 6479 8588 6535
rect 8588 6479 8644 6535
rect 8644 6479 8648 6535
rect 8584 6475 8648 6479
rect 8664 6535 8728 6539
rect 8664 6479 8668 6535
rect 8668 6479 8724 6535
rect 8724 6479 8728 6535
rect 8664 6475 8728 6479
rect 9090 6535 9154 6539
rect 9090 6479 9094 6535
rect 9094 6479 9150 6535
rect 9150 6479 9154 6535
rect 9090 6475 9154 6479
rect 9170 6535 9234 6539
rect 9170 6479 9174 6535
rect 9174 6479 9230 6535
rect 9230 6479 9234 6535
rect 9170 6475 9234 6479
rect 9250 6535 9314 6539
rect 9250 6479 9254 6535
rect 9254 6479 9310 6535
rect 9310 6479 9314 6535
rect 9250 6475 9314 6479
rect 9330 6535 9394 6539
rect 9330 6479 9334 6535
rect 9334 6479 9390 6535
rect 9390 6479 9394 6535
rect 9330 6475 9394 6479
<< metal4 >>
rect 1699 18471 2699 27739
rect 3723 18701 4343 27739
rect 3723 18637 3734 18701
rect 3798 18637 3814 18701
rect 3878 18637 3894 18701
rect 3958 18637 3974 18701
rect 4038 18637 4100 18701
rect 4164 18637 4180 18701
rect 4244 18637 4260 18701
rect 4324 18637 4343 18701
rect 3723 18582 4343 18637
rect 3723 18518 3734 18582
rect 3798 18518 3814 18582
rect 3878 18518 3894 18582
rect 3958 18518 3974 18582
rect 4038 18518 4100 18582
rect 4164 18518 4180 18582
rect 4244 18518 4260 18582
rect 4324 18518 4343 18582
rect 3723 18506 4343 18518
rect 6453 18701 7073 27739
rect 6453 18637 6464 18701
rect 6528 18637 6544 18701
rect 6608 18637 6624 18701
rect 6688 18637 6704 18701
rect 6768 18637 6830 18701
rect 6894 18637 6910 18701
rect 6974 18637 6990 18701
rect 7054 18637 7073 18701
rect 6453 18582 7073 18637
rect 6453 18518 6464 18582
rect 6528 18518 6544 18582
rect 6608 18518 6624 18582
rect 6688 18518 6704 18582
rect 6768 18518 6830 18582
rect 6894 18518 6910 18582
rect 6974 18518 6990 18582
rect 7054 18518 7073 18582
rect 6453 18506 7073 18518
rect 1699 18407 1710 18471
rect 1774 18407 1790 18471
rect 1854 18407 1870 18471
rect 1934 18407 1950 18471
rect 2014 18407 2376 18471
rect 2440 18407 2456 18471
rect 2520 18407 2536 18471
rect 2600 18407 2616 18471
rect 2680 18407 2699 18471
rect 1699 18352 2699 18407
rect 1699 18288 1710 18352
rect 1774 18288 1790 18352
rect 1854 18288 1870 18352
rect 1934 18288 1950 18352
rect 2014 18288 2376 18352
rect 2440 18288 2456 18352
rect 2520 18288 2536 18352
rect 2600 18288 2616 18352
rect 2680 18288 2699 18352
rect 1699 6651 2699 18288
rect 1699 6587 1710 6651
rect 1774 6587 1790 6651
rect 1854 6587 1870 6651
rect 1934 6587 1950 6651
rect 2014 6587 2376 6651
rect 2440 6587 2456 6651
rect 2520 6587 2536 6651
rect 2600 6587 2616 6651
rect 2680 6587 2699 6651
rect 1699 6532 2699 6587
rect 1699 6468 1710 6532
rect 1774 6468 1790 6532
rect 1854 6468 1870 6532
rect 1934 6468 1950 6532
rect 2014 6468 2376 6532
rect 2440 6468 2456 6532
rect 2520 6468 2536 6532
rect 2600 6468 2616 6532
rect 2680 6468 2699 6532
rect 1699 0 2699 6468
rect 8413 18498 9413 27739
rect 8413 18434 8424 18498
rect 8488 18434 8504 18498
rect 8568 18434 8584 18498
rect 8648 18434 8664 18498
rect 8728 18434 9090 18498
rect 9154 18434 9170 18498
rect 9234 18434 9250 18498
rect 9314 18434 9330 18498
rect 9394 18434 9413 18498
rect 8413 18379 9413 18434
rect 8413 18315 8424 18379
rect 8488 18315 8504 18379
rect 8568 18315 8584 18379
rect 8648 18315 8664 18379
rect 8728 18315 9090 18379
rect 9154 18315 9170 18379
rect 9234 18315 9250 18379
rect 9314 18315 9330 18379
rect 9394 18315 9413 18379
rect 8413 6658 9413 18315
rect 8413 6594 8424 6658
rect 8488 6594 8504 6658
rect 8568 6594 8584 6658
rect 8648 6594 8664 6658
rect 8728 6594 9090 6658
rect 9154 6594 9170 6658
rect 9234 6594 9250 6658
rect 9314 6594 9330 6658
rect 9394 6594 9413 6658
rect 8413 6539 9413 6594
rect 8413 6475 8424 6539
rect 8488 6475 8504 6539
rect 8568 6475 8584 6539
rect 8648 6475 8664 6539
rect 8728 6475 9090 6539
rect 9154 6475 9170 6539
rect 9234 6475 9250 6539
rect 9314 6475 9330 6539
rect 9394 6475 9413 6539
rect 8413 0 9413 6475
use sky130_ef_ip__rc_osc_500k  sky130_ef_ip__rc_osc_500k_0
timestamp 1528473026
transform 0 -1 10844 1 0 6464
box 0 0 12242 10724
<< labels >>
flabel metal2 s 5289 27403 5401 28843 0 FreeSans 560 90 0 0 dout
port 1 nsew
flabel metal2 s 5933 27403 6045 28843 0 FreeSans 560 90 0 0 ena
port 2 nsew
flabel metal4 s 3723 18506 4343 27739 0 FreeSans 9600 90 0 0 vssd1
port 3 nsew
flabel metal4 s 6453 18506 7073 27739 0 FreeSans 9600 90 0 0 vccd1
port 4 nsew
flabel metal4 s 1699 0 2699 27739 0 FreeSans 9600 90 0 0 vdda1
port 5 nsew
flabel metal4 s 8413 0 9413 27739 0 FreeSans 9600 90 0 0 vssa1
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 10872 27739
<< end >>
